magic
tech sky130A
magscale 1 2
timestamp 1699112996
<< pwell >>
rect -5762 -1682 5762 1682
<< psubdiff >>
rect -5726 1612 -5630 1646
rect 5630 1612 5726 1646
rect -5726 1550 -5692 1612
rect 5692 1550 5726 1612
rect -5726 -1612 -5692 -1550
rect 5692 -1612 5726 -1550
rect -5726 -1646 -5630 -1612
rect 5630 -1646 5726 -1612
<< psubdiffcont >>
rect -5630 1612 5630 1646
rect -5726 -1550 -5692 1550
rect 5692 -1550 5726 1550
rect -5630 -1646 5630 -1612
<< xpolycontact >>
rect -5596 1084 -5526 1516
rect -5596 -1516 -5526 -1084
rect -5430 1084 -5360 1516
rect -5430 -1516 -5360 -1084
rect -5264 1084 -5194 1516
rect -5264 -1516 -5194 -1084
rect -5098 1084 -5028 1516
rect -5098 -1516 -5028 -1084
rect -4932 1084 -4862 1516
rect -4932 -1516 -4862 -1084
rect -4766 1084 -4696 1516
rect -4766 -1516 -4696 -1084
rect -4600 1084 -4530 1516
rect -4600 -1516 -4530 -1084
rect -4434 1084 -4364 1516
rect -4434 -1516 -4364 -1084
rect -4268 1084 -4198 1516
rect -4268 -1516 -4198 -1084
rect -4102 1084 -4032 1516
rect -4102 -1516 -4032 -1084
rect -3936 1084 -3866 1516
rect -3936 -1516 -3866 -1084
rect -3770 1084 -3700 1516
rect -3770 -1516 -3700 -1084
rect -3604 1084 -3534 1516
rect -3604 -1516 -3534 -1084
rect -3438 1084 -3368 1516
rect -3438 -1516 -3368 -1084
rect -3272 1084 -3202 1516
rect -3272 -1516 -3202 -1084
rect -3106 1084 -3036 1516
rect -3106 -1516 -3036 -1084
rect -2940 1084 -2870 1516
rect -2940 -1516 -2870 -1084
rect -2774 1084 -2704 1516
rect -2774 -1516 -2704 -1084
rect -2608 1084 -2538 1516
rect -2608 -1516 -2538 -1084
rect -2442 1084 -2372 1516
rect -2442 -1516 -2372 -1084
rect -2276 1084 -2206 1516
rect -2276 -1516 -2206 -1084
rect -2110 1084 -2040 1516
rect -2110 -1516 -2040 -1084
rect -1944 1084 -1874 1516
rect -1944 -1516 -1874 -1084
rect -1778 1084 -1708 1516
rect -1778 -1516 -1708 -1084
rect -1612 1084 -1542 1516
rect -1612 -1516 -1542 -1084
rect -1446 1084 -1376 1516
rect -1446 -1516 -1376 -1084
rect -1280 1084 -1210 1516
rect -1280 -1516 -1210 -1084
rect -1114 1084 -1044 1516
rect -1114 -1516 -1044 -1084
rect -948 1084 -878 1516
rect -948 -1516 -878 -1084
rect -782 1084 -712 1516
rect -782 -1516 -712 -1084
rect -616 1084 -546 1516
rect -616 -1516 -546 -1084
rect -450 1084 -380 1516
rect -450 -1516 -380 -1084
rect -284 1084 -214 1516
rect -284 -1516 -214 -1084
rect -118 1084 -48 1516
rect -118 -1516 -48 -1084
rect 48 1084 118 1516
rect 48 -1516 118 -1084
rect 214 1084 284 1516
rect 214 -1516 284 -1084
rect 380 1084 450 1516
rect 380 -1516 450 -1084
rect 546 1084 616 1516
rect 546 -1516 616 -1084
rect 712 1084 782 1516
rect 712 -1516 782 -1084
rect 878 1084 948 1516
rect 878 -1516 948 -1084
rect 1044 1084 1114 1516
rect 1044 -1516 1114 -1084
rect 1210 1084 1280 1516
rect 1210 -1516 1280 -1084
rect 1376 1084 1446 1516
rect 1376 -1516 1446 -1084
rect 1542 1084 1612 1516
rect 1542 -1516 1612 -1084
rect 1708 1084 1778 1516
rect 1708 -1516 1778 -1084
rect 1874 1084 1944 1516
rect 1874 -1516 1944 -1084
rect 2040 1084 2110 1516
rect 2040 -1516 2110 -1084
rect 2206 1084 2276 1516
rect 2206 -1516 2276 -1084
rect 2372 1084 2442 1516
rect 2372 -1516 2442 -1084
rect 2538 1084 2608 1516
rect 2538 -1516 2608 -1084
rect 2704 1084 2774 1516
rect 2704 -1516 2774 -1084
rect 2870 1084 2940 1516
rect 2870 -1516 2940 -1084
rect 3036 1084 3106 1516
rect 3036 -1516 3106 -1084
rect 3202 1084 3272 1516
rect 3202 -1516 3272 -1084
rect 3368 1084 3438 1516
rect 3368 -1516 3438 -1084
rect 3534 1084 3604 1516
rect 3534 -1516 3604 -1084
rect 3700 1084 3770 1516
rect 3700 -1516 3770 -1084
rect 3866 1084 3936 1516
rect 3866 -1516 3936 -1084
rect 4032 1084 4102 1516
rect 4032 -1516 4102 -1084
rect 4198 1084 4268 1516
rect 4198 -1516 4268 -1084
rect 4364 1084 4434 1516
rect 4364 -1516 4434 -1084
rect 4530 1084 4600 1516
rect 4530 -1516 4600 -1084
rect 4696 1084 4766 1516
rect 4696 -1516 4766 -1084
rect 4862 1084 4932 1516
rect 4862 -1516 4932 -1084
rect 5028 1084 5098 1516
rect 5028 -1516 5098 -1084
rect 5194 1084 5264 1516
rect 5194 -1516 5264 -1084
rect 5360 1084 5430 1516
rect 5360 -1516 5430 -1084
rect 5526 1084 5596 1516
rect 5526 -1516 5596 -1084
<< xpolyres >>
rect -5596 -1084 -5526 1084
rect -5430 -1084 -5360 1084
rect -5264 -1084 -5194 1084
rect -5098 -1084 -5028 1084
rect -4932 -1084 -4862 1084
rect -4766 -1084 -4696 1084
rect -4600 -1084 -4530 1084
rect -4434 -1084 -4364 1084
rect -4268 -1084 -4198 1084
rect -4102 -1084 -4032 1084
rect -3936 -1084 -3866 1084
rect -3770 -1084 -3700 1084
rect -3604 -1084 -3534 1084
rect -3438 -1084 -3368 1084
rect -3272 -1084 -3202 1084
rect -3106 -1084 -3036 1084
rect -2940 -1084 -2870 1084
rect -2774 -1084 -2704 1084
rect -2608 -1084 -2538 1084
rect -2442 -1084 -2372 1084
rect -2276 -1084 -2206 1084
rect -2110 -1084 -2040 1084
rect -1944 -1084 -1874 1084
rect -1778 -1084 -1708 1084
rect -1612 -1084 -1542 1084
rect -1446 -1084 -1376 1084
rect -1280 -1084 -1210 1084
rect -1114 -1084 -1044 1084
rect -948 -1084 -878 1084
rect -782 -1084 -712 1084
rect -616 -1084 -546 1084
rect -450 -1084 -380 1084
rect -284 -1084 -214 1084
rect -118 -1084 -48 1084
rect 48 -1084 118 1084
rect 214 -1084 284 1084
rect 380 -1084 450 1084
rect 546 -1084 616 1084
rect 712 -1084 782 1084
rect 878 -1084 948 1084
rect 1044 -1084 1114 1084
rect 1210 -1084 1280 1084
rect 1376 -1084 1446 1084
rect 1542 -1084 1612 1084
rect 1708 -1084 1778 1084
rect 1874 -1084 1944 1084
rect 2040 -1084 2110 1084
rect 2206 -1084 2276 1084
rect 2372 -1084 2442 1084
rect 2538 -1084 2608 1084
rect 2704 -1084 2774 1084
rect 2870 -1084 2940 1084
rect 3036 -1084 3106 1084
rect 3202 -1084 3272 1084
rect 3368 -1084 3438 1084
rect 3534 -1084 3604 1084
rect 3700 -1084 3770 1084
rect 3866 -1084 3936 1084
rect 4032 -1084 4102 1084
rect 4198 -1084 4268 1084
rect 4364 -1084 4434 1084
rect 4530 -1084 4600 1084
rect 4696 -1084 4766 1084
rect 4862 -1084 4932 1084
rect 5028 -1084 5098 1084
rect 5194 -1084 5264 1084
rect 5360 -1084 5430 1084
rect 5526 -1084 5596 1084
<< locali >>
rect -5726 1612 -5630 1646
rect 5630 1612 5726 1646
rect -5726 1550 -5692 1612
rect 5692 1550 5726 1612
rect -5726 -1612 -5692 -1550
rect 5692 -1612 5726 -1550
rect -5726 -1646 -5630 -1612
rect 5630 -1646 5726 -1612
<< viali >>
rect -5580 1101 -5542 1498
rect -5414 1101 -5376 1498
rect -5248 1101 -5210 1498
rect -5082 1101 -5044 1498
rect -4916 1101 -4878 1498
rect -4750 1101 -4712 1498
rect -4584 1101 -4546 1498
rect -4418 1101 -4380 1498
rect -4252 1101 -4214 1498
rect -4086 1101 -4048 1498
rect -3920 1101 -3882 1498
rect -3754 1101 -3716 1498
rect -3588 1101 -3550 1498
rect -3422 1101 -3384 1498
rect -3256 1101 -3218 1498
rect -3090 1101 -3052 1498
rect -2924 1101 -2886 1498
rect -2758 1101 -2720 1498
rect -2592 1101 -2554 1498
rect -2426 1101 -2388 1498
rect -2260 1101 -2222 1498
rect -2094 1101 -2056 1498
rect -1928 1101 -1890 1498
rect -1762 1101 -1724 1498
rect -1596 1101 -1558 1498
rect -1430 1101 -1392 1498
rect -1264 1101 -1226 1498
rect -1098 1101 -1060 1498
rect -932 1101 -894 1498
rect -766 1101 -728 1498
rect -600 1101 -562 1498
rect -434 1101 -396 1498
rect -268 1101 -230 1498
rect -102 1101 -64 1498
rect 64 1101 102 1498
rect 230 1101 268 1498
rect 396 1101 434 1498
rect 562 1101 600 1498
rect 728 1101 766 1498
rect 894 1101 932 1498
rect 1060 1101 1098 1498
rect 1226 1101 1264 1498
rect 1392 1101 1430 1498
rect 1558 1101 1596 1498
rect 1724 1101 1762 1498
rect 1890 1101 1928 1498
rect 2056 1101 2094 1498
rect 2222 1101 2260 1498
rect 2388 1101 2426 1498
rect 2554 1101 2592 1498
rect 2720 1101 2758 1498
rect 2886 1101 2924 1498
rect 3052 1101 3090 1498
rect 3218 1101 3256 1498
rect 3384 1101 3422 1498
rect 3550 1101 3588 1498
rect 3716 1101 3754 1498
rect 3882 1101 3920 1498
rect 4048 1101 4086 1498
rect 4214 1101 4252 1498
rect 4380 1101 4418 1498
rect 4546 1101 4584 1498
rect 4712 1101 4750 1498
rect 4878 1101 4916 1498
rect 5044 1101 5082 1498
rect 5210 1101 5248 1498
rect 5376 1101 5414 1498
rect 5542 1101 5580 1498
rect -5580 -1498 -5542 -1101
rect -5414 -1498 -5376 -1101
rect -5248 -1498 -5210 -1101
rect -5082 -1498 -5044 -1101
rect -4916 -1498 -4878 -1101
rect -4750 -1498 -4712 -1101
rect -4584 -1498 -4546 -1101
rect -4418 -1498 -4380 -1101
rect -4252 -1498 -4214 -1101
rect -4086 -1498 -4048 -1101
rect -3920 -1498 -3882 -1101
rect -3754 -1498 -3716 -1101
rect -3588 -1498 -3550 -1101
rect -3422 -1498 -3384 -1101
rect -3256 -1498 -3218 -1101
rect -3090 -1498 -3052 -1101
rect -2924 -1498 -2886 -1101
rect -2758 -1498 -2720 -1101
rect -2592 -1498 -2554 -1101
rect -2426 -1498 -2388 -1101
rect -2260 -1498 -2222 -1101
rect -2094 -1498 -2056 -1101
rect -1928 -1498 -1890 -1101
rect -1762 -1498 -1724 -1101
rect -1596 -1498 -1558 -1101
rect -1430 -1498 -1392 -1101
rect -1264 -1498 -1226 -1101
rect -1098 -1498 -1060 -1101
rect -932 -1498 -894 -1101
rect -766 -1498 -728 -1101
rect -600 -1498 -562 -1101
rect -434 -1498 -396 -1101
rect -268 -1498 -230 -1101
rect -102 -1498 -64 -1101
rect 64 -1498 102 -1101
rect 230 -1498 268 -1101
rect 396 -1498 434 -1101
rect 562 -1498 600 -1101
rect 728 -1498 766 -1101
rect 894 -1498 932 -1101
rect 1060 -1498 1098 -1101
rect 1226 -1498 1264 -1101
rect 1392 -1498 1430 -1101
rect 1558 -1498 1596 -1101
rect 1724 -1498 1762 -1101
rect 1890 -1498 1928 -1101
rect 2056 -1498 2094 -1101
rect 2222 -1498 2260 -1101
rect 2388 -1498 2426 -1101
rect 2554 -1498 2592 -1101
rect 2720 -1498 2758 -1101
rect 2886 -1498 2924 -1101
rect 3052 -1498 3090 -1101
rect 3218 -1498 3256 -1101
rect 3384 -1498 3422 -1101
rect 3550 -1498 3588 -1101
rect 3716 -1498 3754 -1101
rect 3882 -1498 3920 -1101
rect 4048 -1498 4086 -1101
rect 4214 -1498 4252 -1101
rect 4380 -1498 4418 -1101
rect 4546 -1498 4584 -1101
rect 4712 -1498 4750 -1101
rect 4878 -1498 4916 -1101
rect 5044 -1498 5082 -1101
rect 5210 -1498 5248 -1101
rect 5376 -1498 5414 -1101
rect 5542 -1498 5580 -1101
<< metal1 >>
rect -5586 1498 -5536 1510
rect -5586 1101 -5580 1498
rect -5542 1101 -5536 1498
rect -5586 1089 -5536 1101
rect -5420 1498 -5370 1510
rect -5420 1101 -5414 1498
rect -5376 1101 -5370 1498
rect -5420 1089 -5370 1101
rect -5254 1498 -5204 1510
rect -5254 1101 -5248 1498
rect -5210 1101 -5204 1498
rect -5254 1089 -5204 1101
rect -5088 1498 -5038 1510
rect -5088 1101 -5082 1498
rect -5044 1101 -5038 1498
rect -5088 1089 -5038 1101
rect -4922 1498 -4872 1510
rect -4922 1101 -4916 1498
rect -4878 1101 -4872 1498
rect -4922 1089 -4872 1101
rect -4756 1498 -4706 1510
rect -4756 1101 -4750 1498
rect -4712 1101 -4706 1498
rect -4756 1089 -4706 1101
rect -4590 1498 -4540 1510
rect -4590 1101 -4584 1498
rect -4546 1101 -4540 1498
rect -4590 1089 -4540 1101
rect -4424 1498 -4374 1510
rect -4424 1101 -4418 1498
rect -4380 1101 -4374 1498
rect -4424 1089 -4374 1101
rect -4258 1498 -4208 1510
rect -4258 1101 -4252 1498
rect -4214 1101 -4208 1498
rect -4258 1089 -4208 1101
rect -4092 1498 -4042 1510
rect -4092 1101 -4086 1498
rect -4048 1101 -4042 1498
rect -4092 1089 -4042 1101
rect -3926 1498 -3876 1510
rect -3926 1101 -3920 1498
rect -3882 1101 -3876 1498
rect -3926 1089 -3876 1101
rect -3760 1498 -3710 1510
rect -3760 1101 -3754 1498
rect -3716 1101 -3710 1498
rect -3760 1089 -3710 1101
rect -3594 1498 -3544 1510
rect -3594 1101 -3588 1498
rect -3550 1101 -3544 1498
rect -3594 1089 -3544 1101
rect -3428 1498 -3378 1510
rect -3428 1101 -3422 1498
rect -3384 1101 -3378 1498
rect -3428 1089 -3378 1101
rect -3262 1498 -3212 1510
rect -3262 1101 -3256 1498
rect -3218 1101 -3212 1498
rect -3262 1089 -3212 1101
rect -3096 1498 -3046 1510
rect -3096 1101 -3090 1498
rect -3052 1101 -3046 1498
rect -3096 1089 -3046 1101
rect -2930 1498 -2880 1510
rect -2930 1101 -2924 1498
rect -2886 1101 -2880 1498
rect -2930 1089 -2880 1101
rect -2764 1498 -2714 1510
rect -2764 1101 -2758 1498
rect -2720 1101 -2714 1498
rect -2764 1089 -2714 1101
rect -2598 1498 -2548 1510
rect -2598 1101 -2592 1498
rect -2554 1101 -2548 1498
rect -2598 1089 -2548 1101
rect -2432 1498 -2382 1510
rect -2432 1101 -2426 1498
rect -2388 1101 -2382 1498
rect -2432 1089 -2382 1101
rect -2266 1498 -2216 1510
rect -2266 1101 -2260 1498
rect -2222 1101 -2216 1498
rect -2266 1089 -2216 1101
rect -2100 1498 -2050 1510
rect -2100 1101 -2094 1498
rect -2056 1101 -2050 1498
rect -2100 1089 -2050 1101
rect -1934 1498 -1884 1510
rect -1934 1101 -1928 1498
rect -1890 1101 -1884 1498
rect -1934 1089 -1884 1101
rect -1768 1498 -1718 1510
rect -1768 1101 -1762 1498
rect -1724 1101 -1718 1498
rect -1768 1089 -1718 1101
rect -1602 1498 -1552 1510
rect -1602 1101 -1596 1498
rect -1558 1101 -1552 1498
rect -1602 1089 -1552 1101
rect -1436 1498 -1386 1510
rect -1436 1101 -1430 1498
rect -1392 1101 -1386 1498
rect -1436 1089 -1386 1101
rect -1270 1498 -1220 1510
rect -1270 1101 -1264 1498
rect -1226 1101 -1220 1498
rect -1270 1089 -1220 1101
rect -1104 1498 -1054 1510
rect -1104 1101 -1098 1498
rect -1060 1101 -1054 1498
rect -1104 1089 -1054 1101
rect -938 1498 -888 1510
rect -938 1101 -932 1498
rect -894 1101 -888 1498
rect -938 1089 -888 1101
rect -772 1498 -722 1510
rect -772 1101 -766 1498
rect -728 1101 -722 1498
rect -772 1089 -722 1101
rect -606 1498 -556 1510
rect -606 1101 -600 1498
rect -562 1101 -556 1498
rect -606 1089 -556 1101
rect -440 1498 -390 1510
rect -440 1101 -434 1498
rect -396 1101 -390 1498
rect -440 1089 -390 1101
rect -274 1498 -224 1510
rect -274 1101 -268 1498
rect -230 1101 -224 1498
rect -274 1089 -224 1101
rect -108 1498 -58 1510
rect -108 1101 -102 1498
rect -64 1101 -58 1498
rect -108 1089 -58 1101
rect 58 1498 108 1510
rect 58 1101 64 1498
rect 102 1101 108 1498
rect 58 1089 108 1101
rect 224 1498 274 1510
rect 224 1101 230 1498
rect 268 1101 274 1498
rect 224 1089 274 1101
rect 390 1498 440 1510
rect 390 1101 396 1498
rect 434 1101 440 1498
rect 390 1089 440 1101
rect 556 1498 606 1510
rect 556 1101 562 1498
rect 600 1101 606 1498
rect 556 1089 606 1101
rect 722 1498 772 1510
rect 722 1101 728 1498
rect 766 1101 772 1498
rect 722 1089 772 1101
rect 888 1498 938 1510
rect 888 1101 894 1498
rect 932 1101 938 1498
rect 888 1089 938 1101
rect 1054 1498 1104 1510
rect 1054 1101 1060 1498
rect 1098 1101 1104 1498
rect 1054 1089 1104 1101
rect 1220 1498 1270 1510
rect 1220 1101 1226 1498
rect 1264 1101 1270 1498
rect 1220 1089 1270 1101
rect 1386 1498 1436 1510
rect 1386 1101 1392 1498
rect 1430 1101 1436 1498
rect 1386 1089 1436 1101
rect 1552 1498 1602 1510
rect 1552 1101 1558 1498
rect 1596 1101 1602 1498
rect 1552 1089 1602 1101
rect 1718 1498 1768 1510
rect 1718 1101 1724 1498
rect 1762 1101 1768 1498
rect 1718 1089 1768 1101
rect 1884 1498 1934 1510
rect 1884 1101 1890 1498
rect 1928 1101 1934 1498
rect 1884 1089 1934 1101
rect 2050 1498 2100 1510
rect 2050 1101 2056 1498
rect 2094 1101 2100 1498
rect 2050 1089 2100 1101
rect 2216 1498 2266 1510
rect 2216 1101 2222 1498
rect 2260 1101 2266 1498
rect 2216 1089 2266 1101
rect 2382 1498 2432 1510
rect 2382 1101 2388 1498
rect 2426 1101 2432 1498
rect 2382 1089 2432 1101
rect 2548 1498 2598 1510
rect 2548 1101 2554 1498
rect 2592 1101 2598 1498
rect 2548 1089 2598 1101
rect 2714 1498 2764 1510
rect 2714 1101 2720 1498
rect 2758 1101 2764 1498
rect 2714 1089 2764 1101
rect 2880 1498 2930 1510
rect 2880 1101 2886 1498
rect 2924 1101 2930 1498
rect 2880 1089 2930 1101
rect 3046 1498 3096 1510
rect 3046 1101 3052 1498
rect 3090 1101 3096 1498
rect 3046 1089 3096 1101
rect 3212 1498 3262 1510
rect 3212 1101 3218 1498
rect 3256 1101 3262 1498
rect 3212 1089 3262 1101
rect 3378 1498 3428 1510
rect 3378 1101 3384 1498
rect 3422 1101 3428 1498
rect 3378 1089 3428 1101
rect 3544 1498 3594 1510
rect 3544 1101 3550 1498
rect 3588 1101 3594 1498
rect 3544 1089 3594 1101
rect 3710 1498 3760 1510
rect 3710 1101 3716 1498
rect 3754 1101 3760 1498
rect 3710 1089 3760 1101
rect 3876 1498 3926 1510
rect 3876 1101 3882 1498
rect 3920 1101 3926 1498
rect 3876 1089 3926 1101
rect 4042 1498 4092 1510
rect 4042 1101 4048 1498
rect 4086 1101 4092 1498
rect 4042 1089 4092 1101
rect 4208 1498 4258 1510
rect 4208 1101 4214 1498
rect 4252 1101 4258 1498
rect 4208 1089 4258 1101
rect 4374 1498 4424 1510
rect 4374 1101 4380 1498
rect 4418 1101 4424 1498
rect 4374 1089 4424 1101
rect 4540 1498 4590 1510
rect 4540 1101 4546 1498
rect 4584 1101 4590 1498
rect 4540 1089 4590 1101
rect 4706 1498 4756 1510
rect 4706 1101 4712 1498
rect 4750 1101 4756 1498
rect 4706 1089 4756 1101
rect 4872 1498 4922 1510
rect 4872 1101 4878 1498
rect 4916 1101 4922 1498
rect 4872 1089 4922 1101
rect 5038 1498 5088 1510
rect 5038 1101 5044 1498
rect 5082 1101 5088 1498
rect 5038 1089 5088 1101
rect 5204 1498 5254 1510
rect 5204 1101 5210 1498
rect 5248 1101 5254 1498
rect 5204 1089 5254 1101
rect 5370 1498 5420 1510
rect 5370 1101 5376 1498
rect 5414 1101 5420 1498
rect 5370 1089 5420 1101
rect 5536 1498 5586 1510
rect 5536 1101 5542 1498
rect 5580 1101 5586 1498
rect 5536 1089 5586 1101
rect -5586 -1101 -5536 -1089
rect -5586 -1498 -5580 -1101
rect -5542 -1498 -5536 -1101
rect -5586 -1510 -5536 -1498
rect -5420 -1101 -5370 -1089
rect -5420 -1498 -5414 -1101
rect -5376 -1498 -5370 -1101
rect -5420 -1510 -5370 -1498
rect -5254 -1101 -5204 -1089
rect -5254 -1498 -5248 -1101
rect -5210 -1498 -5204 -1101
rect -5254 -1510 -5204 -1498
rect -5088 -1101 -5038 -1089
rect -5088 -1498 -5082 -1101
rect -5044 -1498 -5038 -1101
rect -5088 -1510 -5038 -1498
rect -4922 -1101 -4872 -1089
rect -4922 -1498 -4916 -1101
rect -4878 -1498 -4872 -1101
rect -4922 -1510 -4872 -1498
rect -4756 -1101 -4706 -1089
rect -4756 -1498 -4750 -1101
rect -4712 -1498 -4706 -1101
rect -4756 -1510 -4706 -1498
rect -4590 -1101 -4540 -1089
rect -4590 -1498 -4584 -1101
rect -4546 -1498 -4540 -1101
rect -4590 -1510 -4540 -1498
rect -4424 -1101 -4374 -1089
rect -4424 -1498 -4418 -1101
rect -4380 -1498 -4374 -1101
rect -4424 -1510 -4374 -1498
rect -4258 -1101 -4208 -1089
rect -4258 -1498 -4252 -1101
rect -4214 -1498 -4208 -1101
rect -4258 -1510 -4208 -1498
rect -4092 -1101 -4042 -1089
rect -4092 -1498 -4086 -1101
rect -4048 -1498 -4042 -1101
rect -4092 -1510 -4042 -1498
rect -3926 -1101 -3876 -1089
rect -3926 -1498 -3920 -1101
rect -3882 -1498 -3876 -1101
rect -3926 -1510 -3876 -1498
rect -3760 -1101 -3710 -1089
rect -3760 -1498 -3754 -1101
rect -3716 -1498 -3710 -1101
rect -3760 -1510 -3710 -1498
rect -3594 -1101 -3544 -1089
rect -3594 -1498 -3588 -1101
rect -3550 -1498 -3544 -1101
rect -3594 -1510 -3544 -1498
rect -3428 -1101 -3378 -1089
rect -3428 -1498 -3422 -1101
rect -3384 -1498 -3378 -1101
rect -3428 -1510 -3378 -1498
rect -3262 -1101 -3212 -1089
rect -3262 -1498 -3256 -1101
rect -3218 -1498 -3212 -1101
rect -3262 -1510 -3212 -1498
rect -3096 -1101 -3046 -1089
rect -3096 -1498 -3090 -1101
rect -3052 -1498 -3046 -1101
rect -3096 -1510 -3046 -1498
rect -2930 -1101 -2880 -1089
rect -2930 -1498 -2924 -1101
rect -2886 -1498 -2880 -1101
rect -2930 -1510 -2880 -1498
rect -2764 -1101 -2714 -1089
rect -2764 -1498 -2758 -1101
rect -2720 -1498 -2714 -1101
rect -2764 -1510 -2714 -1498
rect -2598 -1101 -2548 -1089
rect -2598 -1498 -2592 -1101
rect -2554 -1498 -2548 -1101
rect -2598 -1510 -2548 -1498
rect -2432 -1101 -2382 -1089
rect -2432 -1498 -2426 -1101
rect -2388 -1498 -2382 -1101
rect -2432 -1510 -2382 -1498
rect -2266 -1101 -2216 -1089
rect -2266 -1498 -2260 -1101
rect -2222 -1498 -2216 -1101
rect -2266 -1510 -2216 -1498
rect -2100 -1101 -2050 -1089
rect -2100 -1498 -2094 -1101
rect -2056 -1498 -2050 -1101
rect -2100 -1510 -2050 -1498
rect -1934 -1101 -1884 -1089
rect -1934 -1498 -1928 -1101
rect -1890 -1498 -1884 -1101
rect -1934 -1510 -1884 -1498
rect -1768 -1101 -1718 -1089
rect -1768 -1498 -1762 -1101
rect -1724 -1498 -1718 -1101
rect -1768 -1510 -1718 -1498
rect -1602 -1101 -1552 -1089
rect -1602 -1498 -1596 -1101
rect -1558 -1498 -1552 -1101
rect -1602 -1510 -1552 -1498
rect -1436 -1101 -1386 -1089
rect -1436 -1498 -1430 -1101
rect -1392 -1498 -1386 -1101
rect -1436 -1510 -1386 -1498
rect -1270 -1101 -1220 -1089
rect -1270 -1498 -1264 -1101
rect -1226 -1498 -1220 -1101
rect -1270 -1510 -1220 -1498
rect -1104 -1101 -1054 -1089
rect -1104 -1498 -1098 -1101
rect -1060 -1498 -1054 -1101
rect -1104 -1510 -1054 -1498
rect -938 -1101 -888 -1089
rect -938 -1498 -932 -1101
rect -894 -1498 -888 -1101
rect -938 -1510 -888 -1498
rect -772 -1101 -722 -1089
rect -772 -1498 -766 -1101
rect -728 -1498 -722 -1101
rect -772 -1510 -722 -1498
rect -606 -1101 -556 -1089
rect -606 -1498 -600 -1101
rect -562 -1498 -556 -1101
rect -606 -1510 -556 -1498
rect -440 -1101 -390 -1089
rect -440 -1498 -434 -1101
rect -396 -1498 -390 -1101
rect -440 -1510 -390 -1498
rect -274 -1101 -224 -1089
rect -274 -1498 -268 -1101
rect -230 -1498 -224 -1101
rect -274 -1510 -224 -1498
rect -108 -1101 -58 -1089
rect -108 -1498 -102 -1101
rect -64 -1498 -58 -1101
rect -108 -1510 -58 -1498
rect 58 -1101 108 -1089
rect 58 -1498 64 -1101
rect 102 -1498 108 -1101
rect 58 -1510 108 -1498
rect 224 -1101 274 -1089
rect 224 -1498 230 -1101
rect 268 -1498 274 -1101
rect 224 -1510 274 -1498
rect 390 -1101 440 -1089
rect 390 -1498 396 -1101
rect 434 -1498 440 -1101
rect 390 -1510 440 -1498
rect 556 -1101 606 -1089
rect 556 -1498 562 -1101
rect 600 -1498 606 -1101
rect 556 -1510 606 -1498
rect 722 -1101 772 -1089
rect 722 -1498 728 -1101
rect 766 -1498 772 -1101
rect 722 -1510 772 -1498
rect 888 -1101 938 -1089
rect 888 -1498 894 -1101
rect 932 -1498 938 -1101
rect 888 -1510 938 -1498
rect 1054 -1101 1104 -1089
rect 1054 -1498 1060 -1101
rect 1098 -1498 1104 -1101
rect 1054 -1510 1104 -1498
rect 1220 -1101 1270 -1089
rect 1220 -1498 1226 -1101
rect 1264 -1498 1270 -1101
rect 1220 -1510 1270 -1498
rect 1386 -1101 1436 -1089
rect 1386 -1498 1392 -1101
rect 1430 -1498 1436 -1101
rect 1386 -1510 1436 -1498
rect 1552 -1101 1602 -1089
rect 1552 -1498 1558 -1101
rect 1596 -1498 1602 -1101
rect 1552 -1510 1602 -1498
rect 1718 -1101 1768 -1089
rect 1718 -1498 1724 -1101
rect 1762 -1498 1768 -1101
rect 1718 -1510 1768 -1498
rect 1884 -1101 1934 -1089
rect 1884 -1498 1890 -1101
rect 1928 -1498 1934 -1101
rect 1884 -1510 1934 -1498
rect 2050 -1101 2100 -1089
rect 2050 -1498 2056 -1101
rect 2094 -1498 2100 -1101
rect 2050 -1510 2100 -1498
rect 2216 -1101 2266 -1089
rect 2216 -1498 2222 -1101
rect 2260 -1498 2266 -1101
rect 2216 -1510 2266 -1498
rect 2382 -1101 2432 -1089
rect 2382 -1498 2388 -1101
rect 2426 -1498 2432 -1101
rect 2382 -1510 2432 -1498
rect 2548 -1101 2598 -1089
rect 2548 -1498 2554 -1101
rect 2592 -1498 2598 -1101
rect 2548 -1510 2598 -1498
rect 2714 -1101 2764 -1089
rect 2714 -1498 2720 -1101
rect 2758 -1498 2764 -1101
rect 2714 -1510 2764 -1498
rect 2880 -1101 2930 -1089
rect 2880 -1498 2886 -1101
rect 2924 -1498 2930 -1101
rect 2880 -1510 2930 -1498
rect 3046 -1101 3096 -1089
rect 3046 -1498 3052 -1101
rect 3090 -1498 3096 -1101
rect 3046 -1510 3096 -1498
rect 3212 -1101 3262 -1089
rect 3212 -1498 3218 -1101
rect 3256 -1498 3262 -1101
rect 3212 -1510 3262 -1498
rect 3378 -1101 3428 -1089
rect 3378 -1498 3384 -1101
rect 3422 -1498 3428 -1101
rect 3378 -1510 3428 -1498
rect 3544 -1101 3594 -1089
rect 3544 -1498 3550 -1101
rect 3588 -1498 3594 -1101
rect 3544 -1510 3594 -1498
rect 3710 -1101 3760 -1089
rect 3710 -1498 3716 -1101
rect 3754 -1498 3760 -1101
rect 3710 -1510 3760 -1498
rect 3876 -1101 3926 -1089
rect 3876 -1498 3882 -1101
rect 3920 -1498 3926 -1101
rect 3876 -1510 3926 -1498
rect 4042 -1101 4092 -1089
rect 4042 -1498 4048 -1101
rect 4086 -1498 4092 -1101
rect 4042 -1510 4092 -1498
rect 4208 -1101 4258 -1089
rect 4208 -1498 4214 -1101
rect 4252 -1498 4258 -1101
rect 4208 -1510 4258 -1498
rect 4374 -1101 4424 -1089
rect 4374 -1498 4380 -1101
rect 4418 -1498 4424 -1101
rect 4374 -1510 4424 -1498
rect 4540 -1101 4590 -1089
rect 4540 -1498 4546 -1101
rect 4584 -1498 4590 -1101
rect 4540 -1510 4590 -1498
rect 4706 -1101 4756 -1089
rect 4706 -1498 4712 -1101
rect 4750 -1498 4756 -1101
rect 4706 -1510 4756 -1498
rect 4872 -1101 4922 -1089
rect 4872 -1498 4878 -1101
rect 4916 -1498 4922 -1101
rect 4872 -1510 4922 -1498
rect 5038 -1101 5088 -1089
rect 5038 -1498 5044 -1101
rect 5082 -1498 5088 -1101
rect 5038 -1510 5088 -1498
rect 5204 -1101 5254 -1089
rect 5204 -1498 5210 -1101
rect 5248 -1498 5254 -1101
rect 5204 -1510 5254 -1498
rect 5370 -1101 5420 -1089
rect 5370 -1498 5376 -1101
rect 5414 -1498 5420 -1101
rect 5370 -1510 5420 -1498
rect 5536 -1101 5586 -1089
rect 5536 -1498 5542 -1101
rect 5580 -1498 5586 -1101
rect 5536 -1510 5586 -1498
<< properties >>
string FIXED_BBOX -5709 -1629 5709 1629
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 11 m 1 nx 68 wmin 0.350 lmin 0.50 rho 2000 val 63.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
