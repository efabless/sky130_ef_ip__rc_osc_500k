magic
tech sky130A
timestamp 1699065673
<< pwell >>
rect -139 -150 139 150
<< mvnmos >>
rect -25 -21 25 21
<< mvndiff >>
rect -54 15 -25 21
rect -54 -15 -48 15
rect -31 -15 -25 15
rect -54 -21 -25 -15
rect 25 15 54 21
rect 25 -15 31 15
rect 48 -15 54 15
rect 25 -21 54 -15
<< mvndiffc >>
rect -48 -15 -31 15
rect 31 -15 48 15
<< mvpsubdiff >>
rect -121 126 121 132
rect -121 109 -67 126
rect 67 109 121 126
rect -121 103 121 109
rect -121 78 -92 103
rect -121 -78 -115 78
rect -98 -78 -92 78
rect 92 78 121 103
rect -121 -103 -92 -78
rect 92 -78 98 78
rect 115 -78 121 78
rect 92 -103 121 -78
rect -121 -109 121 -103
rect -121 -126 -67 -109
rect 67 -126 121 -109
rect -121 -132 121 -126
<< mvpsubdiffcont >>
rect -67 109 67 126
rect -115 -78 -98 78
rect 98 -78 115 78
rect -67 -126 67 -109
<< poly >>
rect -25 57 25 65
rect -25 40 -17 57
rect 17 40 25 57
rect -25 21 25 40
rect -25 -40 25 -21
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect -25 -65 25 -57
<< polycont >>
rect -17 40 17 57
rect -17 -57 17 -40
<< locali >>
rect -115 109 -67 126
rect 67 109 115 126
rect -115 78 -98 109
rect 98 78 115 109
rect -25 40 -17 57
rect 17 40 25 57
rect -48 15 -31 23
rect -48 -23 -31 -15
rect 31 15 48 23
rect 31 -23 48 -15
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect -115 -109 -98 -78
rect 98 -109 115 -78
rect -115 -126 -67 -109
rect 67 -126 115 -109
<< viali >>
rect -17 40 17 57
rect -48 -15 -31 15
rect 31 -15 48 15
rect -17 -57 17 -40
<< metal1 >>
rect -23 57 23 60
rect -23 40 -17 57
rect 17 40 23 57
rect -23 37 23 40
rect -51 15 -28 21
rect -51 -15 -48 15
rect -31 -15 -28 15
rect -51 -21 -28 -15
rect 28 15 51 21
rect 28 -15 31 15
rect 48 -15 51 15
rect 28 -21 51 -15
rect -23 -40 23 -37
rect -23 -57 -17 -40
rect 17 -57 23 -40
rect -23 -60 23 -57
<< properties >>
string FIXED_BBOX -106 -117 106 117
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
