magic
tech sky130A
magscale 1 2
timestamp 1699112996
<< metal3 >>
rect -486 612 486 640
rect -486 -612 402 612
rect 466 -612 486 612
rect -486 -640 486 -612
<< via3 >>
rect 402 -612 466 612
<< mimcap >>
rect -446 560 154 600
rect -446 -560 -406 560
rect 114 -560 154 560
rect -446 -600 154 -560
<< mimcapcontact >>
rect -406 -560 114 560
<< metal4 >>
rect 386 612 482 628
rect -407 560 115 561
rect -407 -560 -406 560
rect 114 -560 115 560
rect -407 -561 115 -560
rect 386 -612 402 612
rect 466 -612 482 612
rect 386 -628 482 -612
<< properties >>
string FIXED_BBOX -486 -640 194 640
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.0 l 6.0 val 39.42 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
