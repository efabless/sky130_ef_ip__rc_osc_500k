* NGSPICE file created from sky130_ef_ip__rc_osc_500k.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_6XHUDR a_n242_n264# a_50_n42# a_n108_n42# a_n50_n130#
X0 a_50_n42# a_n50_n130# a_n108_n42# a_n242_n264# sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6ELFTH a_50_n42# a_n50_n139# w_n308_n339# a_n108_n42#
X0 a_50_n42# a_n50_n139# a_n108_n42# w_n308_n339# sky130_fd_pr__pfet_g5v0d10v5 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_L7BSKG a_n73_n11# a_n33_n99# a_15_n11# a_n175_n185#
X0 a_15_n11# a_n33_n99# a_n73_n11# a_n175_n185# sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ a_n2110_1084# a_2206_1084# a_1708_n1516#
+ a_4696_1084# a_48_1084# a_n2442_n1516# a_n1612_1084# a_n4600_1084# a_1708_1084#
+ a_3202_n1516# a_n1446_n1516# a_2870_1084# a_712_1084# a_n284_n1516# a_4696_n1516#
+ a_5028_1084# a_n948_1084# a_2206_n1516# a_n1446_1084# a_n4434_1084# a_n616_n1516#
+ a_3202_1084# a_546_1084# a_1210_n1516# a_n3936_1084# a_5194_n1516# a_2704_1084#
+ a_n4766_n1516# a_n4268_1084# a_3036_1084# a_4198_n1516# a_5526_n1516# a_878_n1516#
+ a_n118_n1516# a_n2442_1084# a_n3770_n1516# a_n5430_1084# a_2538_1084# a_1210_1084#
+ a_5526_1084# a_n5264_n1516# a_4530_n1516# a_n2774_n1516# a_n1944_1084# a_n4932_1084#
+ a_n450_1084# a_n4268_n1516# a_3700_1084# a_3534_n1516# a_n1778_n1516# a_n2276_1084#
+ a_5028_n1516# a_n5264_1084# a_1044_1084# a_4032_1084# a_2538_n1516# a_n3272_n1516#
+ a_n1778_1084# a_n4600_n1516# a_n4766_1084# a_n284_1084# a_n948_n1516# a_3534_1084#
+ a_380_n1516# a_878_1084# a_4032_n1516# a_n2276_n1516# a_n3604_n1516# a_n5098_1084#
+ a_n2940_1084# a_1542_n1516# a_712_n1516# a_3036_n1516# a_n2608_n1516# a_n3272_1084#
+ a_3368_1084# a_2040_1084# a_n1280_n1516# a_n118_1084# a_n4102_n1516# a_n2774_1084#
+ a_2040_n1516# a_1542_1084# a_4530_1084# a_n1612_n1516# a_n5596_n1516# a_4862_n1516#
+ a_n450_n1516# a_n3106_n1516# a_1044_n1516# a_n782_1084# a_214_n1516# a_n3106_1084#
+ a_3866_n1516# a_n5596_1084# a_n1280_1084# a_1376_1084# a_4364_1084# a_n2110_n1516#
+ a_n5726_n1646# a_n2608_1084# a_380_1084# a_5360_n1516# a_n3770_1084# a_n4932_n1516#
+ a_3866_1084# a_n1114_n1516# a_2870_n1516# a_n5098_n1516# a_4364_n1516# a_n616_1084#
+ a_n3936_n1516# a_1874_n1516# a_4198_1084# a_3368_n1516# a_n1114_1084# a_n4102_1084#
+ a_48_n1516# a_n5430_n1516# a_2372_1084# a_5360_1084# a_214_1084# a_n2940_n1516#
+ a_n3604_1084# a_n4434_n1516# a_1874_1084# a_2372_n1516# a_3700_n1516# a_4862_1084#
+ a_n1944_n1516# a_n3438_n1516# a_n782_n1516# a_1376_n1516# a_2704_n1516# a_5194_1084#
+ a_546_n1516# a_n3438_1084#
X0 a_878_1084# a_878_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X1 a_4198_1084# a_4198_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X2 a_n3770_1084# a_n3770_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X3 a_n1446_1084# a_n1446_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X4 a_3700_1084# a_3700_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X5 a_n4268_1084# a_n4268_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X6 a_n2110_1084# a_n2110_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X7 a_1874_1084# a_1874_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X8 a_2372_1084# a_2372_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X9 a_2538_1084# a_2538_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X10 a_4696_1084# a_4696_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X11 a_3036_1084# a_3036_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X12 a_5194_1084# a_5194_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X13 a_n1944_1084# a_n1944_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X14 a_n4766_1084# a_n4766_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X15 a_n2608_1084# a_n2608_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X16 a_n2442_1084# a_n2442_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X17 a_214_1084# a_214_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X18 a_n5430_1084# a_n5430_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X19 a_n5264_1084# a_n5264_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X20 a_n3106_1084# a_n3106_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X21 a_2870_1084# a_2870_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X22 a_n1280_1084# a_n1280_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X23 a_1210_1084# a_1210_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X24 a_3534_1084# a_3534_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X25 a_712_1084# a_712_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X26 a_4032_1084# a_4032_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X27 a_n3604_1084# a_n3604_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X28 a_n118_1084# a_n118_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X29 a_n4102_1084# a_n4102_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X30 a_n1778_1084# a_n1778_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X31 a_4530_1084# a_4530_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X32 a_n4600_1084# a_n4600_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X33 a_n2276_1084# a_n2276_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X34 a_n5098_1084# a_n5098_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X35 a_n616_1084# a_n616_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X36 a_1044_1084# a_1044_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X37 a_3368_1084# a_3368_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X38 a_546_1084# a_546_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X39 a_n2940_1084# a_n2940_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X40 a_n2774_1084# a_n2774_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X41 a_380_1084# a_380_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X42 a_n5596_1084# a_n5596_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X43 a_n3438_1084# a_n3438_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X44 a_n3272_1084# a_n3272_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X45 a_n1114_1084# a_n1114_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X46 a_1708_1084# a_1708_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X47 a_1542_1084# a_1542_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X48 a_2206_1084# a_2206_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X49 a_3866_1084# a_3866_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X50 a_2040_1084# a_2040_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X51 a_4364_1084# a_4364_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X52 a_5028_1084# a_5028_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X53 a_n450_1084# a_n450_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X54 a_n3936_1084# a_n3936_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X55 a_n1612_1084# a_n1612_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X56 a_n284_1084# a_n284_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X57 a_n4434_1084# a_n4434_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X58 a_48_1084# a_48_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X59 a_2704_1084# a_2704_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X60 a_4862_1084# a_4862_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X61 a_3202_1084# a_3202_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X62 a_5360_1084# a_5360_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X63 a_5526_1084# a_5526_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X64 a_n948_1084# a_n948_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X65 a_n782_1084# a_n782_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X66 a_n4932_1084# a_n4932_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
X67 a_1376_1084# a_1376_n1516# a_n5726_n1646# sky130_fd_pr__res_xhigh_po_0p35 l=10.8
.ends

.subckt sky130_fd_pr__pfet_01v8_LGS3BL a_n73_n64# a_n33_n161# a_15_n64# w_n211_n284#
X0 a_15_n64# a_n33_n161# a_n73_n64# w_n211_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_64Z3AY a_15_n131# a_n175_n243# a_n33_91# a_n73_n131#
X0 a_15_n131# a_n33_91# a_n73_n131# a_n175_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt level_shifter dvdd out_h outb_h in_l inb_l avss avdd dvss
XXM15 outb_h out_h avdd m1_1336_n1198# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM16 avdd outb_h avdd m1_1336_n1198# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM17 avss outb_h avss in_l sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM18 avss avss out_h inb_l sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM19 m1_2204_n1198# out_h avdd avdd sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM7 dvdd in_l inb_l dvdd sky130_fd_pr__pfet_01v8_LGS3BL
XXM8 inb_l dvss in_l dvss sky130_fd_pr__nfet_01v8_64Z3AY
XXM20 m1_2204_n1198# outb_h avdd out_h sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
.ends

.subckt sky130_fd_pr__nfet_01v8_L9WNCD a_15_n19# a_n175_n193# a_n73_n19# a_n33_n107#
X0 a_15_n19# a_n33_n107# a_n73_n19# a_n175_n193# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ a_n147_n147# a_n45_n45#
D0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_AZFCP3 m3_n486_n640# c1_n446_n600#
X0 c1_n446_n600# m3_n486_n640# sky130_fd_pr__cap_mim_m3_1 l=6 w=3
.ends

.subckt sky130_fd_pr__pfet_01v8_2Z69BZ w_n211_n226# a_n73_n6# a_15_n6# a_n33_n103#
X0 a_15_n6# a_n33_n103# a_n73_n6# w_n211_n226# sky130_fd_pr__pfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt sky130_ef_ip__rc_osc_500k avdd avss dvss dvdd ena dout
XXM12 avss m1_11932_n1089# avss m1_7381_n511# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM34 avdd level_shifter_0/out_h avdd m1_6724_n888# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM23 avss m1_9629_n1544# m1_4901_916# level_shifter_0/out_h sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM35 dout level_shifter_0/inb_l dvss dvss sky130_fd_pr__nfet_01v8_L7BSKG
XXM13 avss m1_12146_n889# m1_11932_n1089# ena sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM25 avdd m1_6724_n888# avdd m1_7989_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM24 avdd m1_6724_n888# avdd m1_7373_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM36 avss m1_6949_n1486# m1_6724_n888# level_shifter_0/out_h sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM37 m1_7381_n511# m1_10298_n888# avdd m1_11069_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM15 m1_9735_n892# m1_9177_n893# avdd m1_9837_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM26 avdd m1_6724_n888# avdd m1_8605_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM38 avss m1_7381_n511# m1_10628_n1035# m1_10298_n888# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM16 avss m1_9735_n892# m1_9516_n1035# m1_9177_n893# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM27 avss m1_8404_n1035# avss m1_9629_n1544# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM39 avdd m1_6724_n888# avdd m1_10453_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM17 avdd m1_6724_n888# avdd m1_9221_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM28 avss m1_7848_n1035# avss m1_9629_n1544# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM18 avdd m1_6724_n888# avdd m1_9837_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM29 avss m1_7292_n1035# avss m1_9629_n1544# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM19 avss m1_9516_n1035# avss m1_9629_n1544# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
Xsky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_0 m1_8408_n2556# m1_12724_n2556# m1_12226_n5156#
+ m1_15048_n2556# m1_10400_n2556# m1_7910_n5156# m1_8740_n2556# m1_5752_n2556# m1_12060_n2556#
+ m1_13554_n5156# m1_8906_n5156# m1_13388_n2556# m1_11064_n2556# m1_10234_n5156# m1_15214_n5156#
+ m1_15380_n2556# m1_9404_n2556# m1_12558_n5156# m1_9072_n2556# m1_6084_n2556# m1_9902_n5156#
+ m1_13720_n2556# m1_11064_n2556# m1_11562_n5156# m1_6416_n2556# m1_15546_n5156# m1_13056_n2556#
+ m1_5586_n5156# m1_6084_n2556# m1_13388_n2556# m1_14550_n5156# m1_15878_n5156# m1_11230_n5156#
+ m1_10234_n5156# m1_8076_n2556# m1_6582_n5156# m1_5088_n2556# m1_13056_n2556# m1_11728_n2556#
+ m1_14882_n1618# m1_5254_n5156# m1_14882_n5156# m1_7578_n5156# m1_8408_n2556# m1_5420_n2556#
+ m1_10068_n2556# m1_6250_n5156# m1_14052_n2556# m1_13886_n5156# m1_8574_n5156# m1_8076_n2556#
+ m1_15546_n5156# m1_5088_n2556# m1_11396_n2556# m1_14384_n2556# m1_12890_n5156# m1_7246_n5156#
+ m1_8740_n2556# m1_5918_n5156# m1_5752_n2556# m1_10068_n2556# m1_9570_n5156# m1_14052_n2556#
+ m1_10898_n5156# m1_11396_n2556# m1_14550_n5156# m1_8242_n5156# m1_6914_n5156# m1_5420_n2556#
+ m1_7412_n2556# m1_11894_n5156# m1_11230_n5156# m1_13554_n5156# m1_7910_n5156# m1_7080_n2556#
+ m1_13720_n2556# m1_12392_n2556# m1_9238_n5156# m1_10400_n2556# m1_6250_n5156# m1_7744_n2556#
+ m1_12558_n5156# m1_12060_n2556# m1_15048_n2556# m1_8906_n5156# m1_4922_n5156# m1_15214_n5156#
+ m1_9902_n5156# m1_7246_n5156# m1_11562_n5156# m1_9736_n2556# m1_10566_n5156# m1_7412_n2556#
+ m1_14218_n5156# avdd m1_9072_n2556# m1_11728_n2556# m1_14716_n2556# m1_8242_n5156#
+ avss m1_7744_n2556# m1_10732_n2556# m1_15878_n5156# m1_6748_n2556# m1_5586_n5156#
+ m1_14384_n2556# m1_9238_n5156# m1_13222_n5156# m1_5254_n5156# m1_14882_n5156# m1_9736_n2556#
+ m1_6582_n5156# m1_12226_n5156# m1_14716_n2556# m1_13886_n5156# m1_9404_n2556# m1_6416_n2556#
+ m1_10566_n5156# m1_4922_n5156# m1_12724_n2556# m1_15712_n2556# m1_10732_n2556# m1_7578_n5156#
+ m1_6748_n2556# m1_5918_n5156# m1_12392_n2556# m1_12890_n5156# m1_14218_n5156# m1_15380_n2556#
+ m1_8574_n5156# m1_6914_n5156# m1_9570_n5156# m1_11894_n5156# m1_13222_n5156# m1_15712_n2556#
+ m1_10898_n5156# m1_7080_n2556# sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ
Xsky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_1 m1_8222_4094# m1_12538_4094# m1_12040_1494#
+ m1_15194_4094# m1_10546_4094# m1_8056_1494# m1_8886_4094# m1_5898_4094# m1_12206_4094#
+ m1_13700_1494# m1_9052_1494# m1_13202_4094# m1_11210_4094# m1_10048_1494# m1_15028_1494#
+ m1_15526_4094# m1_9550_4094# m1_12704_1494# m1_8886_4094# m1_5898_4094# m1_9716_1494#
+ m1_13534_4094# m1_10878_4094# m1_11708_1494# m1_6562_4094# m1_15692_1494# m1_13202_4094#
+ m1_5732_1494# m1_6230_4094# m1_13534_4094# m1_14696_1494# m1_14882_n1618# m1_11376_1494#
+ m1_10380_1494# m1_7890_4094# m1_6728_1494# m1_4902_4094# m1_12870_4094# m1_11542_4094#
+ m1_15858_4094# m1_5068_1494# m1_15028_1494# m1_7724_1494# m1_8554_4094# m1_5566_4094#
+ m1_9882_4094# m1_6064_1494# m1_14198_4094# m1_14032_1494# m1_8720_1494# m1_8222_4094#
+ m1_15360_1494# m1_5234_4094# m1_11542_4094# m1_14530_4094# m1_13036_1494# m1_7060_1494#
+ m1_8554_4094# m1_5732_1494# m1_5566_4094# m1_10214_4094# m1_9384_1494# m1_13866_4094#
+ m1_10712_1494# m1_11210_4094# m1_14364_1494# m1_8056_1494# m1_6728_1494# m1_5234_4094#
+ m1_7558_4094# m1_12040_1494# m1_11044_1494# m1_13368_1494# m1_7724_1494# m1_7226_4094#
+ m1_13866_4094# m1_12538_4094# m1_9052_1494# m1_10214_4094# m1_6396_1494# m1_7558_4094#
+ m1_12372_1494# m1_11874_4094# m1_14862_4094# m1_8720_1494# m1_4901_916# m1_15360_1494#
+ m1_10048_1494# m1_7392_1494# m1_11376_1494# m1_9550_4094# m1_10712_1494# m1_7226_4094#
+ m1_14364_1494# m1_4902_4094# m1_9218_4094# m1_11874_4094# m1_14862_4094# m1_8388_1494#
+ avss m1_7890_4094# m1_10878_4094# m1_15692_1494# m1_6562_4094# m1_5400_1494# m1_14198_4094#
+ m1_9384_1494# m1_13368_1494# m1_5400_1494# m1_14696_1494# m1_9882_4094# m1_6396_1494#
+ m1_12372_1494# m1_14530_4094# m1_13700_1494# m1_9218_4094# m1_6230_4094# m1_10380_1494#
+ m1_5068_1494# m1_12870_4094# m1_15858_4094# m1_10546_4094# m1_7392_1494# m1_6894_4094#
+ m1_6064_1494# m1_12206_4094# m1_12704_1494# m1_14032_1494# m1_15194_4094# m1_8388_1494#
+ m1_7060_1494# m1_9716_1494# m1_11708_1494# m1_13036_1494# m1_15526_4094# m1_11044_1494#
+ m1_6894_4094# sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ
XXM1 avss m1_7516_n887# m1_7292_n1035# m1_7381_n511# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM2 m1_7516_n887# m1_7381_n511# avdd m1_7373_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM3 m1_8067_n893# m1_7516_n887# avdd m1_7989_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
Xlevel_shifter_0 dvdd level_shifter_0/out_h level_shifter_0/outb_h ena level_shifter_0/inb_l
+ avss avdd dvss level_shifter
XXM4 avss m1_8067_n893# m1_7848_n1035# m1_7516_n887# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
Xsky130_fd_pr__nfet_01v8_L9WNCD_0 m1_16326_216# dvss dvss m1_12146_n889# sky130_fd_pr__nfet_01v8_L9WNCD
XXM5 m1_16326_216# dvss dout ena sky130_fd_pr__nfet_01v8_L9WNCD
XD3 dvss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
XXM7 m1_9177_n893# m1_8623_n885# avdd m1_9221_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM9 m1_8623_n885# m1_8067_n893# avdd m1_8605_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM8 avss m1_9177_n893# m1_8960_n1035# m1_8623_n885# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
Xsky130_fd_pr__pfet_01v8_LGS3BL_0 dvdd m1_12146_n889# dout dvdd sky130_fd_pr__pfet_01v8_LGS3BL
XXC1 avss m1_7516_n887# sky130_fd_pr__cap_mim_m3_1_AZFCP3
XXC2 avss m1_8067_n893# sky130_fd_pr__cap_mim_m3_1_AZFCP3
XXC3 avss m1_8623_n885# sky130_fd_pr__cap_mim_m3_1_AZFCP3
XXC4 avss m1_9177_n893# sky130_fd_pr__cap_mim_m3_1_AZFCP3
Xsky130_fd_pr__pfet_01v8_2Z69BZ_0 dvdd m1_12146_n889# dvdd ena sky130_fd_pr__pfet_01v8_2Z69BZ
Xsky130_fd_pr__cap_mim_m3_1_AZFCP3_1 avss m1_9735_n892# sky130_fd_pr__cap_mim_m3_1_AZFCP3
XXM40 avdd m1_6724_n888# avdd m1_11069_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM41 avss m1_10628_n1035# avss m1_9629_n1544# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM30 avss m1_6949_n1486# avss m1_9629_n1544# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM31 m1_10298_n888# m1_9735_n892# avdd m1_10453_n21# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM42 avss m1_10072_n1035# avss m1_9629_n1544# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM20 avss m1_8960_n1035# avss m1_9629_n1544# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM32 avss m1_10298_n888# m1_10072_n1035# m1_9735_n892# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM10 avss m1_8623_n885# m1_8404_n1035# m1_8067_n893# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM21 avss m1_9629_n1544# avss m1_9629_n1544# sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
XXM11 m1_12146_n889# m1_7381_n511# avdd dvdd sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM22 avdd m1_6724_n888# avdd m1_6724_n888# sky130_fd_pr__pfet_g5v0d10v5_6ELFTH
XXM33 avss m1_9629_n1544# avss level_shifter_0/outb_h sky130_fd_pr__nfet_g5v0d10v5_6XHUDR
.ends

