magic
tech sky130A
magscale 1 2
timestamp 1699295625
<< dnwell >>
rect 4504 1092 16514 4934
rect 4504 -1720 14362 1092
rect 4504 -5558 16514 -1720
<< nwell >>
rect 4388 4728 16630 5050
rect 4388 -5352 4710 4728
rect 16308 1298 16630 4728
rect 11506 360 12376 1039
rect 14156 976 16630 1298
rect 11506 -318 11760 360
rect 14156 -1604 14478 976
rect 16001 -633 16055 -281
rect 14156 -1926 16630 -1604
rect 16308 -5352 16630 -1926
rect 4388 -5674 16630 -5352
<< mvnsubdiff >>
rect 4461 4957 16557 4977
rect 4461 4923 4541 4957
rect 16477 4923 16557 4957
rect 4461 4903 16557 4923
rect 4461 4897 4535 4903
rect 4461 -5521 4481 4897
rect 4515 -5521 4535 4897
rect 16483 4897 16557 4903
rect 16483 1143 16503 4897
rect 16537 1143 16557 4897
rect 16483 1123 16557 1143
rect 14331 1103 16557 1123
rect 14331 1069 14436 1103
rect 16467 1069 16557 1103
rect 14331 1049 16557 1069
rect 14331 1021 14405 1049
rect 14331 -1645 14351 1021
rect 14385 -1645 14405 1021
rect 14331 -1677 14405 -1645
rect 14331 -1697 16557 -1677
rect 14331 -1731 14436 -1697
rect 16466 -1731 16557 -1697
rect 14331 -1751 16557 -1731
rect 4461 -5527 4535 -5521
rect 16483 -1765 16557 -1751
rect 16483 -5521 16503 -1765
rect 16537 -5521 16557 -1765
rect 16483 -5527 16557 -5521
rect 4461 -5547 16557 -5527
rect 4461 -5581 4541 -5547
rect 16477 -5581 16557 -5547
rect 4461 -5601 16557 -5581
<< mvnsubdiffcont >>
rect 4541 4923 16477 4957
rect 4481 -5521 4515 4897
rect 16503 1143 16537 4897
rect 14436 1069 16467 1103
rect 14351 -1645 14385 1021
rect 14436 -1731 16466 -1697
rect 16503 -5521 16537 -1765
rect 4541 -5581 16477 -5547
<< locali >>
rect 4474 4957 16539 4962
rect 4474 4923 4541 4957
rect 16477 4923 16539 4957
rect 4474 4897 16539 4923
rect 4474 -5521 4481 4897
rect 4515 4819 16503 4897
rect 4515 2009 4598 4819
rect 4581 -1669 4598 2009
rect 4683 4621 16332 4735
rect 4683 1416 4797 4621
rect 16218 1416 16332 4621
rect 4683 1397 16332 1416
rect 4683 1312 12690 1397
rect 14131 1312 16332 1397
rect 4683 1302 16332 1312
rect 16434 4012 16503 4819
rect 16537 4819 16539 4897
rect 16434 2038 16442 4012
rect 4884 -361 6024 1302
rect 16434 1219 16503 2038
rect 6569 1077 12273 1078
rect 6522 1051 12273 1077
rect 6522 994 6607 1051
rect 12250 994 12273 1051
rect 6522 919 12273 994
rect 6522 476 6676 919
rect 11953 477 12273 919
rect 14243 1192 16503 1219
rect 14243 1167 14419 1192
rect 6522 250 6891 476
rect 7165 250 7507 476
rect 7781 250 8123 476
rect 8397 250 8739 476
rect 9013 250 9355 476
rect 9629 250 9971 476
rect 10245 250 10587 476
rect 10861 250 11203 476
rect 11953 476 12397 477
rect 11477 250 12397 476
rect 6522 -205 6676 250
rect 12269 -205 12397 250
rect 6522 -362 12397 -205
rect 6569 -363 12397 -362
rect 6569 -364 12288 -363
rect 12265 -468 12388 -467
rect 5408 -627 12388 -468
rect 5408 -1063 5539 -627
rect 10979 -1056 11841 -627
rect 5408 -1225 5510 -1063
rect 10979 -1067 11184 -1056
rect 5666 -1069 11184 -1067
rect 5666 -1226 6049 -1069
rect 6304 -1226 6605 -1069
rect 6860 -1226 7161 -1069
rect 7416 -1226 7717 -1069
rect 7972 -1226 8273 -1069
rect 8528 -1226 8829 -1069
rect 9084 -1226 9385 -1069
rect 9640 -1226 9941 -1069
rect 10196 -1226 10497 -1069
rect 10752 -1225 11184 -1069
rect 11340 -1067 11841 -1056
rect 12265 -1067 12388 -627
rect 11340 -1225 12388 -1067
rect 10752 -1226 12388 -1225
rect 12265 -1661 12388 -1226
rect 4515 -5475 4598 -1669
rect 5519 -1711 12388 -1661
rect 5519 -1746 12293 -1711
rect 5519 -1801 5571 -1746
rect 12246 -1801 12293 -1746
rect 14243 -1731 14268 1167
rect 14333 1127 14419 1167
rect 15845 1143 16503 1192
rect 15845 1127 16537 1143
rect 14333 1103 16537 1127
rect 14333 1069 14436 1103
rect 16467 1069 16537 1103
rect 14333 1057 16537 1069
rect 14333 1021 14392 1057
rect 14333 -1645 14351 1021
rect 14385 -1645 14392 1021
rect 14907 899 15312 906
rect 14907 770 15021 899
rect 14907 268 15312 770
rect 15984 576 16437 578
rect 14581 60 15312 268
rect 15979 575 16437 576
rect 15979 448 16011 575
rect 16215 448 16437 575
rect 15979 445 16437 448
rect 15979 349 16122 445
rect 15979 286 16004 349
rect 16111 286 16122 349
rect 15979 123 16122 286
rect 15979 93 16437 123
rect 14840 -183 15312 60
rect 15981 48 16437 93
rect 15981 -134 16437 -59
rect 14576 -198 15312 -183
rect 14576 -199 15201 -198
rect 14576 -426 14619 -199
rect 14792 -426 15201 -199
rect 15983 -278 16126 -134
rect 14576 -440 15201 -426
rect 15960 -286 16126 -278
rect 15960 -482 15989 -286
rect 16123 -482 16126 -286
rect 15960 -543 16126 -482
rect 15960 -617 16442 -543
rect 15964 -618 16442 -617
rect 15645 -848 15965 -717
rect 16012 -735 16442 -660
rect 14605 -989 14811 -987
rect 14605 -991 15978 -989
rect 16012 -991 16127 -735
rect 14605 -1001 16127 -991
rect 14605 -1161 14619 -1001
rect 14796 -1037 16127 -1001
rect 14796 -1161 16442 -1037
rect 14605 -1176 16442 -1161
rect 14333 -1657 14392 -1645
rect 14333 -1697 16537 -1657
rect 14333 -1731 14436 -1697
rect 16466 -1731 16537 -1697
rect 14243 -1765 16537 -1731
rect 14243 -1781 16503 -1765
rect 5519 -1820 12293 -1801
rect 4694 -1903 16339 -1885
rect 4694 -1906 9762 -1903
rect 4694 -1985 6250 -1906
rect 7909 -1982 9762 -1906
rect 11421 -1982 16339 -1903
rect 7909 -1985 16339 -1982
rect 4694 -1999 16339 -1985
rect 4694 -2629 4808 -1999
rect 4694 -4590 4707 -2629
rect 4801 -4590 4808 -2629
rect 4694 -5247 4808 -4590
rect 16225 -2628 16339 -1999
rect 16225 -4589 16228 -2628
rect 16322 -4589 16339 -2628
rect 16225 -5247 16339 -4589
rect 4694 -5361 16339 -5247
rect 16434 -5475 16503 -1781
rect 4515 -5521 16503 -5475
rect 4474 -5547 16537 -5521
rect 4474 -5581 4541 -5547
rect 16477 -5581 16537 -5547
<< viali >>
rect 4500 -1669 4515 2009
rect 4515 -1669 4581 2009
rect 12690 1312 14131 1397
rect 16442 2038 16503 4012
rect 16503 2038 16530 4012
rect 6607 994 12250 1051
rect 12707 873 14111 1206
rect 6891 250 7165 477
rect 7507 250 7781 477
rect 8123 250 8397 477
rect 8739 250 9013 477
rect 9355 250 9629 477
rect 9971 250 10245 477
rect 10587 250 10861 477
rect 11203 250 11477 477
rect 5510 -1232 5666 -1063
rect 6049 -1226 6304 -1069
rect 6605 -1226 6860 -1069
rect 7161 -1226 7416 -1069
rect 7717 -1226 7972 -1069
rect 8273 -1226 8528 -1069
rect 8829 -1226 9084 -1069
rect 9385 -1226 9640 -1069
rect 9941 -1226 10196 -1069
rect 10497 -1226 10752 -1069
rect 11184 -1225 11340 -1056
rect 5571 -1801 12246 -1746
rect 12700 -1751 14104 -1418
rect 14268 -1731 14333 1167
rect 14419 1127 15845 1192
rect 15021 770 15317 899
rect 16011 448 16215 575
rect 16004 286 16111 349
rect 14619 -426 14792 -199
rect 15989 -482 16123 -286
rect 14619 -1161 14796 -1001
rect 6250 -1985 7909 -1906
rect 9762 -1982 11421 -1903
rect 4707 -4590 4801 -2629
rect 16228 -4589 16322 -2628
<< metal1 >>
rect 4902 4094 5138 4526
rect 5234 4094 5470 4526
rect 5566 4094 5802 4526
rect 5898 4094 6134 4526
rect 6230 4094 6466 4526
rect 6562 4094 6798 4526
rect 6894 4094 7130 4526
rect 7226 4094 7462 4526
rect 7558 4094 7794 4526
rect 7890 4094 8126 4526
rect 8222 4094 8458 4526
rect 8554 4094 8790 4526
rect 8886 4094 9122 4526
rect 9218 4094 9454 4526
rect 9550 4094 9786 4526
rect 9882 4094 10118 4526
rect 10214 4094 10450 4526
rect 10546 4094 10782 4526
rect 10878 4094 11114 4526
rect 11210 4094 11446 4526
rect 11542 4094 11778 4526
rect 11874 4094 12110 4526
rect 12206 4094 12442 4526
rect 12538 4094 12774 4526
rect 12870 4094 13106 4526
rect 13202 4094 13438 4526
rect 13534 4094 13770 4526
rect 13866 4094 14102 4526
rect 14198 4094 14434 4526
rect 14530 4094 14766 4526
rect 14862 4094 15098 4526
rect 15194 4094 15430 4526
rect 15526 4094 15762 4526
rect 15858 4094 16094 4526
rect 16436 4012 16536 4024
rect 16432 2038 16442 4012
rect 16530 2038 16540 4012
rect 16436 2026 16536 2038
rect 4494 2009 4587 2021
rect 4490 -1669 4500 2009
rect 4581 789 4591 2009
rect 4901 967 4976 1927
rect 5068 1494 5304 1926
rect 5400 1494 5636 1926
rect 5732 1494 5968 1926
rect 6064 1494 6300 1926
rect 6396 1494 6632 1926
rect 6728 1494 6964 1926
rect 7060 1494 7296 1926
rect 7392 1494 7628 1926
rect 7724 1494 7960 1926
rect 8056 1494 8292 1926
rect 8388 1494 8624 1926
rect 8720 1494 8956 1926
rect 9052 1494 9288 1926
rect 9384 1494 9620 1926
rect 9716 1494 9952 1926
rect 10048 1494 10284 1926
rect 10380 1494 10616 1926
rect 10712 1494 10948 1926
rect 11044 1494 11280 1926
rect 11376 1494 11612 1926
rect 11708 1494 11944 1926
rect 12040 1494 12276 1926
rect 12372 1494 12608 1926
rect 12704 1494 12940 1926
rect 13036 1494 13272 1926
rect 13368 1494 13604 1926
rect 13700 1494 13936 1926
rect 14032 1494 14268 1926
rect 14364 1494 14600 1926
rect 14696 1494 14932 1926
rect 15028 1494 15264 1926
rect 15360 1494 15596 1926
rect 15692 1494 15928 1926
rect 5015 1406 6216 1409
rect 12673 1406 14156 1416
rect 5015 1397 14156 1406
rect 5015 1395 12690 1397
rect 5015 1268 5042 1395
rect 6183 1312 12690 1395
rect 14131 1312 14156 1397
rect 6183 1268 14156 1312
rect 5015 1251 14156 1268
rect 5195 1250 14156 1251
rect 12673 1227 14156 1250
rect 14225 1325 15882 1350
rect 14225 1227 14265 1325
rect 15846 1227 15882 1325
rect 12673 1206 14155 1227
rect 6525 1144 12301 1174
rect 6525 1079 6578 1144
rect 12274 1079 12301 1144
rect 6525 1051 12301 1079
rect 6525 994 6607 1051
rect 12250 994 12301 1051
rect 6525 984 12301 994
rect 4901 916 6227 967
rect 4581 -364 6020 789
rect 4581 -1669 4591 -364
rect 5827 -728 5837 -707
rect 5582 -1051 5666 -803
rect 5736 -954 5764 -737
rect 5772 -768 5837 -728
rect 5827 -769 5837 -768
rect 5994 -769 6004 -707
rect 5504 -1063 5672 -1051
rect 5500 -1232 5510 -1063
rect 5666 -1232 5676 -1063
rect 5504 -1244 5672 -1232
rect 5842 -1545 5874 -806
rect 6176 -884 6227 916
rect 12673 873 12707 1206
rect 14111 873 14155 1206
rect 6761 801 11250 848
rect 12673 832 14155 873
rect 14225 1192 15882 1227
rect 14225 1167 14419 1192
rect 6761 22 6808 801
rect 6871 591 6902 801
rect 6961 483 7061 741
rect 6879 477 7177 483
rect 6879 250 6891 477
rect 7165 250 7177 477
rect 6879 244 7177 250
rect 6724 -25 6808 22
rect 6348 -611 6358 -590
rect 6291 -652 6358 -611
rect 6515 -611 6525 -590
rect 6515 -648 6605 -611
rect 6515 -652 6525 -648
rect 6291 -952 6328 -652
rect 6037 -1069 6316 -1063
rect 6037 -1226 6049 -1069
rect 6304 -1226 6316 -1069
rect 6037 -1232 6316 -1226
rect 6135 -1489 6219 -1232
rect 6292 -1545 6325 -1346
rect 6397 -1545 6437 -795
rect 6568 -922 6605 -648
rect 6724 -888 6771 -25
rect 6870 -586 6902 128
rect 6976 -22 7080 244
rect 7373 -21 7417 748
rect 7487 591 7518 801
rect 7577 483 7677 741
rect 7495 477 7793 483
rect 7495 250 7507 477
rect 7781 250 7793 477
rect 7495 244 7793 250
rect 7480 -346 7519 133
rect 7381 -511 7391 -346
rect 7448 -388 7519 -346
rect 7578 -158 7617 60
rect 7989 -21 8033 748
rect 8103 591 8134 801
rect 8193 483 8293 741
rect 8111 477 8409 483
rect 8111 250 8123 477
rect 8397 250 8409 477
rect 8111 244 8409 250
rect 7578 -248 7592 -158
rect 7802 -248 7812 -158
rect 7578 -348 7617 -248
rect 8096 -348 8135 133
rect 7578 -387 8135 -348
rect 8207 -158 8246 64
rect 8605 -21 8649 748
rect 8719 591 8750 801
rect 8809 483 8909 741
rect 8727 477 9025 483
rect 8727 250 8739 477
rect 9013 250 9025 477
rect 8727 244 9025 250
rect 8207 -248 8223 -158
rect 8433 -248 8443 -158
rect 8207 -346 8246 -248
rect 8712 -346 8751 133
rect 8207 -385 8751 -346
rect 8833 -158 8872 71
rect 9221 -21 9265 748
rect 9335 591 9366 801
rect 9425 483 9525 741
rect 9343 477 9641 483
rect 9343 250 9355 477
rect 9629 250 9641 477
rect 9343 244 9641 250
rect 8833 -248 8855 -158
rect 9065 -248 9075 -158
rect 8833 -346 8872 -248
rect 9328 -346 9367 133
rect 8833 -385 9367 -346
rect 9436 -158 9475 63
rect 9837 -21 9881 748
rect 9951 591 9982 801
rect 10041 483 10141 741
rect 9959 477 10257 483
rect 9959 250 9971 477
rect 10245 250 10257 477
rect 9959 244 10257 250
rect 9436 -248 9459 -158
rect 9669 -248 9679 -158
rect 9436 -346 9475 -248
rect 9944 -346 9983 133
rect 9436 -385 9983 -346
rect 10060 -176 10099 70
rect 10453 -21 10497 748
rect 10567 591 10598 801
rect 10657 483 10757 741
rect 10575 477 10873 483
rect 10575 250 10587 477
rect 10861 250 10873 477
rect 10575 244 10873 250
rect 10262 -176 10272 -158
rect 10060 -232 10272 -176
rect 10060 -346 10099 -232
rect 10262 -248 10272 -232
rect 10482 -248 10492 -158
rect 10560 -346 10599 133
rect 10060 -385 10599 -346
rect 10671 -346 10710 67
rect 11069 -21 11113 748
rect 11183 591 11214 801
rect 11273 483 11373 741
rect 11890 499 11900 598
rect 12260 499 12270 598
rect 11191 477 11489 483
rect 11191 250 11203 477
rect 11477 250 11489 477
rect 11191 244 11489 250
rect 11176 -346 11215 133
rect 11293 -342 11332 70
rect 11899 -8 11983 499
rect 12408 293 12418 314
rect 12146 255 12418 293
rect 12044 -161 12088 150
rect 11591 -205 12088 -161
rect 10671 -385 11215 -346
rect 7448 -511 7458 -388
rect 6860 -648 6870 -586
rect 7027 -648 7037 -586
rect 6847 -922 6884 -715
rect 6568 -959 6884 -922
rect 6593 -1069 6872 -1063
rect 6593 -1226 6605 -1069
rect 6860 -1226 6872 -1069
rect 6593 -1232 6872 -1226
rect 6691 -1243 6783 -1232
rect 6699 -1486 6783 -1243
rect 6849 -1544 6882 -1341
rect 6949 -1486 6991 -797
rect 7292 -993 7334 -800
rect 7404 -954 7443 -511
rect 7578 -659 7617 -387
rect 7516 -698 7617 -659
rect 7516 -887 7555 -698
rect 7848 -993 7890 -800
rect 7960 -954 7999 -387
rect 8207 -658 8246 -385
rect 8067 -697 8246 -658
rect 8067 -893 8106 -697
rect 8404 -993 8446 -800
rect 8516 -954 8555 -385
rect 8833 -656 8872 -385
rect 8623 -695 8872 -656
rect 8623 -885 8662 -695
rect 8960 -993 9002 -800
rect 9072 -954 9111 -385
rect 9436 -653 9475 -385
rect 9177 -692 9475 -653
rect 9177 -893 9216 -692
rect 9516 -993 9558 -800
rect 9628 -954 9667 -385
rect 10060 -654 10099 -385
rect 9735 -693 10099 -654
rect 9735 -892 9774 -693
rect 10072 -993 10114 -800
rect 10184 -954 10223 -385
rect 10671 -647 10710 -385
rect 10298 -686 10710 -647
rect 10298 -888 10337 -686
rect 10628 -993 10670 -800
rect 10740 -954 10779 -385
rect 11280 -507 11290 -342
rect 11347 -384 11357 -342
rect 11591 -384 11635 -205
rect 11347 -451 11635 -384
rect 11347 -507 11357 -451
rect 11293 -642 11332 -507
rect 10845 -681 11332 -642
rect 10845 -887 10884 -681
rect 7292 -1035 7547 -993
rect 7848 -1035 8103 -993
rect 8404 -1035 8659 -993
rect 8960 -1035 9215 -993
rect 9516 -1035 9771 -993
rect 10072 -1035 10327 -993
rect 10628 -1035 10883 -993
rect 7149 -1069 7428 -1063
rect 7149 -1226 7161 -1069
rect 7416 -1226 7428 -1069
rect 7149 -1232 7428 -1226
rect 7247 -1243 7339 -1232
rect 7255 -1486 7339 -1243
rect 7405 -1544 7438 -1341
rect 7505 -1486 7547 -1035
rect 7705 -1069 7984 -1063
rect 7705 -1226 7717 -1069
rect 7972 -1226 7984 -1069
rect 7705 -1232 7984 -1226
rect 7803 -1243 7895 -1232
rect 7811 -1486 7895 -1243
rect 7961 -1544 7994 -1341
rect 8061 -1486 8103 -1035
rect 8261 -1069 8540 -1063
rect 8261 -1226 8273 -1069
rect 8528 -1226 8540 -1069
rect 8261 -1232 8540 -1226
rect 8359 -1243 8451 -1232
rect 8367 -1486 8451 -1243
rect 8517 -1544 8550 -1341
rect 8617 -1486 8659 -1035
rect 8817 -1069 9096 -1063
rect 8817 -1226 8829 -1069
rect 9084 -1226 9096 -1069
rect 8817 -1232 9096 -1226
rect 8915 -1243 9007 -1232
rect 8923 -1486 9007 -1243
rect 9073 -1544 9106 -1341
rect 9173 -1486 9215 -1035
rect 9373 -1069 9652 -1063
rect 9373 -1226 9385 -1069
rect 9640 -1226 9652 -1069
rect 9373 -1232 9652 -1226
rect 9471 -1243 9563 -1232
rect 9479 -1486 9563 -1243
rect 9629 -1544 9662 -1341
rect 9729 -1486 9771 -1035
rect 9929 -1069 10208 -1063
rect 9929 -1226 9941 -1069
rect 10196 -1226 10208 -1069
rect 9929 -1232 10208 -1226
rect 10027 -1243 10119 -1232
rect 10035 -1486 10119 -1243
rect 10185 -1544 10218 -1341
rect 10285 -1486 10327 -1035
rect 10485 -1069 10764 -1063
rect 10485 -1226 10497 -1069
rect 10752 -1226 10764 -1069
rect 10485 -1232 10764 -1226
rect 10583 -1243 10675 -1232
rect 10591 -1486 10675 -1243
rect 10741 -1544 10774 -1341
rect 10841 -1486 10883 -1035
rect 11178 -1056 11346 -1044
rect 11178 -1061 11184 -1056
rect 11044 -1069 11184 -1061
rect 11044 -1226 11053 -1069
rect 11340 -1225 11346 -1056
rect 11308 -1226 11346 -1225
rect 11044 -1235 11346 -1226
rect 11178 -1237 11346 -1235
rect 11591 -1227 11635 -451
rect 11932 -1051 11970 -814
rect 12037 -931 12073 -741
rect 12146 -889 12184 255
rect 12408 236 12418 255
rect 12609 236 12619 314
rect 12438 -529 12717 -495
rect 12438 -713 12472 -529
rect 12318 -777 12328 -713
rect 12515 -777 12525 -713
rect 12037 -967 12457 -931
rect 12421 -1036 12457 -967
rect 11932 -1089 12183 -1051
rect 12421 -1075 12485 -1036
rect 11212 -1400 11296 -1237
rect 11591 -1270 12078 -1227
rect 11649 -1271 12078 -1270
rect 11212 -1401 11972 -1400
rect 11212 -1483 11982 -1401
rect 11212 -1484 11870 -1483
rect 5842 -1593 10792 -1545
rect 12034 -1550 12078 -1271
rect 12145 -1484 12183 -1089
rect 12475 -1100 12485 -1075
rect 12672 -1100 12682 -1036
rect 14225 -1358 14268 1167
rect 14113 -1368 14268 -1358
rect 12656 -1418 14268 -1368
rect 4494 -1681 4587 -1669
rect 5517 -1746 12291 -1661
rect 5517 -1801 5571 -1746
rect 12246 -1801 12291 -1746
rect 12656 -1751 12700 -1418
rect 14104 -1731 14268 -1418
rect 14333 1127 14419 1167
rect 15845 1127 15882 1192
rect 14333 1100 15882 1127
rect 14333 -1731 14402 1100
rect 16046 1028 16121 1933
rect 14882 953 16121 1028
rect 14655 809 14665 881
rect 14841 809 14851 881
rect 14642 314 14695 514
rect 14779 428 14841 809
rect 14453 242 14463 314
rect 14639 260 14695 314
rect 14639 242 14649 260
rect 14740 106 14772 390
rect 14628 34 14638 106
rect 14814 34 14824 106
rect 14740 -33 14772 -31
rect 14600 -105 14610 -33
rect 14786 -105 14796 -33
rect 14605 -199 14811 -181
rect 14605 -426 14619 -199
rect 14792 -426 14811 -199
rect 14605 -1001 14811 -426
rect 14605 -1161 14619 -1001
rect 14796 -1161 14811 -1001
rect 14605 -1174 14811 -1161
rect 14882 -1543 14957 953
rect 15009 899 15329 905
rect 15009 770 15021 899
rect 15317 770 15329 899
rect 16252 890 16630 1447
rect 15009 764 15329 770
rect 15530 880 16630 890
rect 15530 781 15541 880
rect 15901 781 16630 880
rect 15530 690 16630 781
rect 15026 503 15036 602
rect 15396 503 15406 602
rect 15530 575 16227 690
rect 15032 -740 15194 503
rect 15530 448 16011 575
rect 16215 448 16227 575
rect 15530 442 16227 448
rect 15530 365 16017 442
rect 15530 349 16226 365
rect 15530 286 16004 349
rect 16111 286 16226 349
rect 15530 271 16226 286
rect 15530 269 15730 271
rect 16217 270 16226 271
rect 16326 264 16374 370
rect 16326 216 16448 264
rect 16206 155 16292 209
rect 15877 -19 15887 -2
rect 15816 -74 15887 -19
rect 16063 -11 16073 -2
rect 16206 -11 16247 155
rect 16063 -60 16247 -11
rect 16063 -74 16073 -60
rect 15816 -384 15854 -74
rect 16206 -243 16247 -60
rect 16275 -61 16285 108
rect 16354 -61 16364 108
rect 16298 -144 16364 -61
rect 15983 -286 16129 -274
rect 15726 -422 15854 -384
rect 15726 -538 15764 -422
rect 15891 -452 15989 -286
rect 15823 -482 15989 -452
rect 16123 -482 16229 -286
rect 15823 -484 16229 -482
rect 15823 -494 16129 -484
rect 15823 -534 16103 -494
rect 15641 -648 15651 -576
rect 15827 -648 15837 -576
rect 15891 -740 16103 -534
rect 16323 -547 16364 -144
rect 15032 -940 16103 -740
rect 16175 -588 16364 -547
rect 16175 -888 16216 -588
rect 16400 -636 16448 216
rect 16327 -684 16448 -636
rect 16327 -888 16375 -684
rect 15543 -1283 16103 -940
rect 16165 -1003 16175 -944
rect 16361 -1003 16371 -944
rect 15543 -1483 16630 -1283
rect 14882 -1618 16121 -1543
rect 14104 -1751 14402 -1731
rect 12656 -1782 14402 -1751
rect 5517 -1818 12291 -1801
rect 6238 -1906 7921 -1900
rect 6238 -1985 6250 -1906
rect 7909 -1985 7921 -1906
rect 6238 -1991 7921 -1985
rect 9750 -1903 11433 -1897
rect 9750 -1982 9762 -1903
rect 11421 -1982 11433 -1903
rect 9750 -1988 11433 -1982
rect 4474 -2131 4993 -2124
rect 4474 -2540 4488 -2131
rect 4739 -2540 4993 -2131
rect 4474 -2556 4993 -2540
rect 5088 -2556 5324 -2124
rect 5420 -2556 5656 -2124
rect 5752 -2556 5988 -2124
rect 6084 -2556 6320 -2124
rect 6416 -2556 6652 -2124
rect 6748 -2556 6984 -2124
rect 7080 -2556 7316 -2124
rect 7412 -2556 7648 -2124
rect 7744 -2556 7980 -2124
rect 8076 -2556 8312 -2124
rect 8408 -2556 8644 -2124
rect 8740 -2556 8976 -2124
rect 9072 -2556 9308 -2124
rect 9404 -2556 9640 -2124
rect 9736 -2556 9972 -2124
rect 10068 -2556 10304 -2124
rect 10400 -2556 10636 -2124
rect 10732 -2556 10968 -2124
rect 11064 -2556 11300 -2124
rect 11396 -2556 11632 -2124
rect 11728 -2556 11964 -2124
rect 12060 -2556 12296 -2124
rect 12392 -2556 12628 -2124
rect 12724 -2556 12960 -2124
rect 13056 -2556 13292 -2124
rect 13388 -2556 13624 -2124
rect 13720 -2556 13956 -2124
rect 14052 -2556 14288 -2124
rect 14384 -2556 14620 -2124
rect 14716 -2556 14952 -2124
rect 15048 -2556 15284 -2124
rect 15380 -2556 15616 -2124
rect 15712 -2556 15948 -2124
rect 16046 -2559 16121 -1618
rect 16252 -2040 16630 -1483
rect 4701 -2629 4807 -2617
rect 16222 -2628 16328 -2616
rect 4697 -4590 4707 -2629
rect 4801 -4590 4811 -2629
rect 16218 -4589 16228 -2628
rect 16322 -4589 16332 -2628
rect 4701 -4602 4807 -4590
rect 16222 -4601 16328 -4589
rect 4922 -5156 5158 -4724
rect 5254 -5156 5490 -4724
rect 5586 -5156 5822 -4724
rect 5918 -5156 6154 -4724
rect 6250 -5156 6486 -4724
rect 6582 -5156 6818 -4724
rect 6914 -5156 7150 -4724
rect 7246 -5156 7482 -4724
rect 7578 -5156 7814 -4724
rect 7910 -5156 8146 -4724
rect 8242 -5156 8478 -4724
rect 8574 -5156 8810 -4724
rect 8906 -5156 9142 -4724
rect 9238 -5156 9474 -4724
rect 9570 -5156 9806 -4724
rect 9902 -5156 10138 -4724
rect 10234 -5156 10470 -4724
rect 10566 -5156 10802 -4724
rect 10898 -5156 11134 -4724
rect 11230 -5156 11466 -4724
rect 11562 -5156 11798 -4724
rect 11894 -5156 12130 -4724
rect 12226 -5156 12462 -4724
rect 12558 -5156 12794 -4724
rect 12890 -5156 13126 -4724
rect 13222 -5156 13458 -4724
rect 13554 -5156 13790 -4724
rect 13886 -5156 14122 -4724
rect 14218 -5156 14454 -4724
rect 14550 -5156 14786 -4724
rect 14882 -5156 15118 -4724
rect 15214 -5156 15450 -4724
rect 15546 -5156 15782 -4724
rect 15878 -5156 16114 -4724
<< via1 >>
rect 16442 2038 16530 4012
rect 4500 -1669 4581 2009
rect 5042 1268 6183 1395
rect 14265 1227 15846 1325
rect 6578 1079 12274 1144
rect 5837 -769 5994 -707
rect 5510 -1232 5666 -1063
rect 12707 873 14111 1206
rect 6891 250 7165 477
rect 6358 -652 6515 -590
rect 6049 -1226 6304 -1069
rect 7507 250 7781 477
rect 7391 -511 7448 -346
rect 8123 250 8397 477
rect 7592 -248 7802 -158
rect 8739 250 9013 477
rect 8223 -248 8433 -158
rect 9355 250 9629 477
rect 8855 -248 9065 -158
rect 9971 250 10245 477
rect 9459 -248 9669 -158
rect 10587 250 10861 477
rect 10272 -248 10482 -158
rect 11900 499 12260 598
rect 11203 250 11477 477
rect 6870 -648 7027 -586
rect 6605 -1226 6860 -1069
rect 11290 -507 11347 -342
rect 7161 -1226 7416 -1069
rect 7717 -1226 7972 -1069
rect 8273 -1226 8528 -1069
rect 8829 -1226 9084 -1069
rect 9385 -1226 9640 -1069
rect 9941 -1226 10196 -1069
rect 10497 -1226 10752 -1069
rect 11053 -1225 11184 -1069
rect 11184 -1225 11308 -1069
rect 11053 -1226 11308 -1225
rect 12418 236 12609 314
rect 12328 -777 12515 -713
rect 12485 -1100 12672 -1036
rect 5571 -1801 12246 -1746
rect 12700 -1751 14104 -1418
rect 14665 809 14841 881
rect 14463 242 14639 314
rect 14638 34 14814 106
rect 14610 -105 14786 -33
rect 15021 770 15317 899
rect 15541 781 15901 880
rect 15036 503 15396 602
rect 15887 -74 16063 -2
rect 16285 -61 16354 108
rect 15651 -648 15827 -576
rect 16175 -1003 16361 -944
rect 6250 -1985 7909 -1906
rect 9762 -1982 11421 -1903
rect 4488 -2540 4739 -2131
rect 4707 -4590 4801 -2629
rect 16228 -4589 16322 -2628
<< metal2 >>
rect 16442 4021 16530 4022
rect 4388 4012 16630 4021
rect 4388 2038 16442 4012
rect 16530 2038 16630 4012
rect 4388 2027 16630 2038
rect 4480 2009 4746 2027
rect 4480 -1669 4500 2009
rect 4581 -1669 4746 2009
rect 5015 1395 6216 1409
rect 5015 1391 5042 1395
rect 4480 -2131 4746 -1669
rect 4480 -2540 4488 -2131
rect 4739 -2540 4746 -2131
rect 4480 -2546 4746 -2540
rect 5013 1268 5042 1391
rect 6183 1268 6216 1395
rect 5013 1251 6216 1268
rect 5013 790 5563 1251
rect 6841 1191 8499 2027
rect 9797 1191 11455 2027
rect 12673 1227 14156 1416
rect 14225 1325 15882 2027
rect 14225 1227 14265 1325
rect 15846 1227 15882 1325
rect 12673 1206 14155 1227
rect 14225 1208 15882 1227
rect 6507 1144 12342 1191
rect 6507 1079 6578 1144
rect 12274 1079 12342 1144
rect 6507 981 12342 1079
rect 5013 -367 6023 790
rect 6841 525 8499 981
rect 9797 525 11455 981
rect 12673 873 12707 1206
rect 14111 873 14155 1206
rect 15021 900 15317 909
rect 12673 832 14155 873
rect 14651 899 15906 900
rect 14651 881 15021 899
rect 14651 809 14665 881
rect 14841 809 15021 881
rect 14651 770 15021 809
rect 15317 880 15906 899
rect 15317 781 15541 880
rect 15901 781 15906 880
rect 15317 770 15906 781
rect 14651 768 15906 770
rect 15021 760 15317 768
rect 11900 600 12260 608
rect 15036 602 15396 612
rect 11900 598 15036 600
rect 6519 477 11554 525
rect 12260 503 15036 598
rect 12260 502 15396 503
rect 11900 489 12260 499
rect 15036 493 15396 502
rect 6519 250 6891 477
rect 7165 250 7507 477
rect 7781 250 8123 477
rect 8397 250 8739 477
rect 9013 250 9355 477
rect 9629 250 9971 477
rect 10245 250 10587 477
rect 10861 250 11203 477
rect 11477 250 11554 477
rect 6519 209 11554 250
rect 12418 314 12609 324
rect 14463 314 14639 324
rect 12609 255 14360 299
rect 14462 255 14463 299
rect 12418 226 12609 236
rect 14316 202 14360 255
rect 14639 255 15962 299
rect 14463 232 14639 242
rect 14316 158 15812 202
rect 14638 106 14814 116
rect 14638 24 14814 34
rect 15768 -20 15812 158
rect 15918 85 15962 255
rect 16285 108 16354 118
rect 15918 41 16285 85
rect 15887 -2 16063 8
rect 14610 -33 14786 -23
rect 6909 -82 7007 -72
rect 7975 -82 8073 -72
rect 7592 -151 7802 -148
rect 7007 -158 7802 -151
rect 7007 -248 7592 -158
rect 7007 -256 7802 -248
rect 7592 -258 7802 -256
rect 6909 -307 7007 -297
rect 9041 -82 9139 -72
rect 8073 -148 8239 -147
rect 8073 -158 8433 -148
rect 8073 -248 8223 -158
rect 8073 -257 8433 -248
rect 8223 -258 8433 -257
rect 8855 -158 9041 -148
rect 10107 -82 10205 -72
rect 8855 -258 9041 -248
rect 7975 -307 8073 -297
rect 9459 -158 10107 -148
rect 9669 -248 10107 -158
rect 9459 -257 10107 -248
rect 9459 -258 9669 -257
rect 9041 -307 9139 -297
rect 11173 -82 11271 -72
rect 10470 -148 11173 -147
rect 10272 -158 11173 -148
rect 10482 -248 11173 -158
rect 10272 -257 11173 -248
rect 10272 -258 10482 -257
rect 10107 -307 10205 -297
rect 11173 -307 11271 -297
rect 7391 -346 7448 -336
rect 5013 -1030 5563 -367
rect 11290 -342 11347 -332
rect 7448 -454 11290 -413
rect 7391 -521 7448 -511
rect 11290 -517 11347 -507
rect 6358 -590 6515 -580
rect 6870 -586 7027 -576
rect 6320 -651 6358 -590
rect 6515 -648 6870 -590
rect 7027 -648 12651 -590
rect 6515 -651 12651 -648
rect 6358 -662 6515 -652
rect 6870 -658 7027 -651
rect 5837 -707 5994 -697
rect 12318 -713 12515 -703
rect 12318 -724 12328 -713
rect 5994 -769 12328 -724
rect 5837 -779 5994 -769
rect 12328 -787 12515 -777
rect 12590 -748 12651 -651
rect 12590 -809 12926 -748
rect 5013 -1063 11523 -1030
rect 12485 -1035 12672 -1026
rect 14076 -1035 14141 -74
rect 15768 -64 15887 -20
rect 16430 85 16630 156
rect 16354 41 16630 85
rect 16430 -44 16630 41
rect 16285 -71 16354 -61
rect 15887 -84 16063 -74
rect 14610 -115 14786 -105
rect 15404 -283 15957 -229
rect 15651 -576 15827 -566
rect 15903 -588 15957 -283
rect 15827 -635 15957 -588
rect 15651 -658 15827 -648
rect 15903 -761 15957 -635
rect 16430 -761 16630 -688
rect 15903 -815 16630 -761
rect 16242 -934 16298 -815
rect 16430 -888 16630 -815
rect 16175 -944 16361 -934
rect 16175 -1013 16361 -1003
rect 5013 -1232 5510 -1063
rect 5666 -1069 11523 -1063
rect 5666 -1226 6049 -1069
rect 6304 -1226 6605 -1069
rect 6860 -1226 7161 -1069
rect 7416 -1226 7717 -1069
rect 7972 -1226 8273 -1069
rect 8528 -1226 8829 -1069
rect 9084 -1226 9385 -1069
rect 9640 -1226 9941 -1069
rect 10196 -1226 10497 -1069
rect 10752 -1226 11053 -1069
rect 11308 -1226 11523 -1069
rect 12483 -1036 14141 -1035
rect 12483 -1100 12485 -1036
rect 12672 -1100 14141 -1036
rect 12485 -1110 12672 -1100
rect 5666 -1232 11523 -1226
rect 5013 -1332 11523 -1232
rect 5013 -1636 5563 -1332
rect 6249 -1636 7908 -1332
rect 9763 -1636 11422 -1332
rect 12656 -1418 14138 -1368
rect 5013 -1746 12318 -1636
rect 5013 -1801 5571 -1746
rect 12246 -1801 12318 -1746
rect 12656 -1751 12700 -1418
rect 14104 -1751 14138 -1418
rect 12656 -1782 14138 -1751
rect 5013 -1850 12318 -1801
rect 5013 -2612 5563 -1850
rect 6249 -1906 7909 -1850
rect 6249 -1985 6250 -1906
rect 6249 -1995 7909 -1985
rect 9762 -1903 11422 -1850
rect 11421 -1982 11422 -1903
rect 9762 -1992 11422 -1982
rect 6249 -2612 7908 -1995
rect 9763 -2612 11422 -1992
rect 4388 -2628 16630 -2612
rect 4388 -2629 16228 -2628
rect 4388 -4590 4707 -2629
rect 4801 -2666 16228 -2629
rect 4801 -2933 7479 -2666
rect 11865 -2933 16228 -2666
rect 4801 -4589 16228 -2933
rect 16322 -4589 16630 -2628
rect 4801 -4590 16630 -4589
rect 4388 -4606 16630 -4590
<< via2 >>
rect 6909 -297 7007 -82
rect 7975 -297 8073 -82
rect 9041 -158 9139 -82
rect 9041 -248 9065 -158
rect 9065 -248 9139 -158
rect 9041 -297 9139 -248
rect 10107 -297 10205 -82
rect 11173 -297 11271 -82
rect 7479 -2933 11865 -2666
<< metal3 >>
rect 6899 -82 7017 -77
rect 6899 -297 6909 -82
rect 7007 -297 7017 -82
rect 6899 -302 7017 -297
rect 7965 -82 8083 -77
rect 7965 -297 7975 -82
rect 8073 -297 8083 -82
rect 7965 -302 8083 -297
rect 9031 -82 9149 -77
rect 9031 -297 9041 -82
rect 9139 -297 9149 -82
rect 9031 -302 9149 -297
rect 10097 -82 10215 -77
rect 10097 -297 10107 -82
rect 10205 -297 10215 -82
rect 10097 -302 10215 -297
rect 11163 -82 11281 -77
rect 11163 -297 11173 -82
rect 11271 -297 11281 -82
rect 11163 -302 11281 -297
rect 7592 -1744 7686 -464
rect 8658 -1744 8752 -464
rect 9724 -1743 9818 -463
rect 10790 -1743 10884 -463
rect 7482 -2103 7492 -1853
rect 7590 -2103 7600 -1853
rect 7482 -2661 7600 -2103
rect 8548 -2103 8558 -1853
rect 8656 -2103 8666 -1853
rect 8548 -2661 8666 -2103
rect 9614 -2103 9624 -1853
rect 9722 -2103 9732 -1853
rect 9614 -2661 9732 -2103
rect 10680 -2103 10690 -1853
rect 10788 -2103 10798 -1853
rect 10680 -2661 10798 -2103
rect 11746 -2103 11756 -1853
rect 11854 -2103 11864 -1853
rect 11746 -2661 11864 -2103
rect 7469 -2666 11875 -2661
rect 7469 -2933 7479 -2666
rect 11865 -2933 11875 -2666
rect 7469 -2938 11875 -2933
<< via3 >>
rect 6909 -297 7007 -82
rect 7975 -297 8073 -82
rect 9041 -297 9139 -82
rect 10107 -297 10205 -82
rect 11173 -297 11271 -82
rect 7492 -2103 7590 -1853
rect 8558 -2103 8656 -1853
rect 9624 -2103 9722 -1853
rect 10690 -2103 10788 -1853
rect 11756 -2103 11854 -1853
<< metal4 >>
rect 6898 -82 7018 -76
rect 6898 -297 6909 -82
rect 7007 -297 7018 -82
rect 6898 -304 7018 -297
rect 7964 -82 8084 -76
rect 7964 -297 7975 -82
rect 8073 -297 8084 -82
rect 7964 -304 8084 -297
rect 9030 -82 9150 -76
rect 9030 -297 9041 -82
rect 9139 -297 9150 -82
rect 9030 -304 9150 -297
rect 10096 -82 10216 -76
rect 10096 -297 10107 -82
rect 10205 -297 10216 -82
rect 10096 -304 10216 -297
rect 11162 -82 11282 -76
rect 11162 -297 11173 -82
rect 11271 -297 11282 -82
rect 11162 -304 11282 -297
rect 6909 -1346 7007 -304
rect 7975 -1346 8073 -304
rect 9041 -1346 9139 -304
rect 10107 -1346 10205 -304
rect 11173 -1346 11271 -304
rect 7492 -1852 7590 -1594
rect 8558 -1852 8656 -1594
rect 9624 -1852 9722 -1594
rect 10690 -1852 10788 -1594
rect 11756 -1852 11854 -1594
rect 7491 -1853 7591 -1852
rect 7491 -2103 7492 -1853
rect 7590 -2103 7591 -1853
rect 7491 -2104 7591 -2103
rect 8557 -1853 8657 -1852
rect 8557 -2103 8558 -1853
rect 8656 -2103 8657 -1853
rect 8557 -2104 8657 -2103
rect 9623 -1853 9723 -1852
rect 9623 -2103 9624 -1853
rect 9722 -2103 9723 -1853
rect 9623 -2104 9723 -2103
rect 10689 -1853 10789 -1852
rect 10689 -2103 10690 -1853
rect 10788 -2103 10789 -1853
rect 10689 -2104 10789 -2103
rect 11755 -1853 11855 -1852
rect 11755 -2103 11756 -1853
rect 11854 -2103 11855 -1853
rect 11755 -2104 11855 -2103
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D3
timestamp 1699295625
transform 1 0 14727 0 1 -70
box -183 -183 183 183
use level_shifter  level_shifter_0
timestamp 1699295625
transform -1 0 15320 0 -1 -1460
box -422 -2544 2736 144
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  sky130_fd_pr__cap_mim_m3_1_AZFCP3_1
timestamp 1699295625
transform 1 0 11370 0 1 -1103
box -486 -640 486 640
use sky130_fd_pr__nfet_01v8_L9WNCD  sky130_fd_pr__nfet_01v8_L9WNCD_0
timestamp 1699295625
transform 1 0 16263 0 1 284
box -211 -229 211 229
use sky130_fd_pr__pfet_01v8_2Z69BZ  sky130_fd_pr__pfet_01v8_2Z69BZ_0
timestamp 1699295625
transform 1 0 15790 0 1 -529
box -211 -226 211 226
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0
timestamp 1699295625
transform 1 0 16266 0 -1 -349
box -211 -284 211 284
use sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ  sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_0
timestamp 1699295625
transform 1 0 10518 0 1 -3640
box -5762 -1682 5762 1682
use sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ  sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_1
timestamp 1699295625
transform 1 0 10498 0 1 3010
box -5762 -1682 5762 1682
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC1
timestamp 1699295625
transform 1 0 7106 0 1 -1104
box -486 -640 486 640
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC2
timestamp 1699295625
transform 1 0 8172 0 1 -1104
box -486 -640 486 640
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC3
timestamp 1699295625
transform 1 0 9238 0 1 -1103
box -486 -640 486 640
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC4
timestamp 1699295625
transform 1 0 10304 0 1 -1103
box -486 -640 486 640
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM1
timestamp 1699295625
transform 1 0 7420 0 1 -844
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM2
timestamp 1699295625
transform 1 0 7502 0 1 21
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM3
timestamp 1699295625
transform 1 0 8118 0 1 21
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM4
timestamp 1699295625
transform 1 0 7976 0 1 -844
box -278 -300 278 300
use sky130_fd_pr__nfet_01v8_L9WNCD  XM5
timestamp 1699295625
transform 1 0 16270 0 1 -880
box -211 -229 211 229
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM7
timestamp 1699295625
transform 1 0 9350 0 1 21
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM8
timestamp 1699295625
transform 1 0 9088 0 1 -844
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM9
timestamp 1699295625
transform 1 0 8734 0 1 21
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM10
timestamp 1699295625
transform 1 0 8532 0 1 -844
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM11
timestamp 1699295625
transform 1 0 12068 0 1 21
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM12
timestamp 1699295625
transform 1 0 12056 0 1 -1446
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM13
timestamp 1699295625
transform 1 0 12056 0 1 -846
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM15
timestamp 1699295625
transform 1 0 9966 0 1 21
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM16
timestamp 1699295625
transform 1 0 9644 0 1 -844
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM17
timestamp 1699295625
transform 1 0 9350 0 1 699
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM18
timestamp 1699295625
transform 1 0 9966 0 1 699
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM19
timestamp 1699295625
transform 1 0 9644 0 1 -1444
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM20
timestamp 1699295625
transform 1 0 9088 0 1 -1444
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM21
timestamp 1699295625
transform 1 0 6308 0 1 -1444
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM22
timestamp 1699295625
transform 1 0 6886 0 1 699
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM23
timestamp 1699295625
transform 1 0 6308 0 1 -846
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM24
timestamp 1699295625
transform 1 0 7502 0 1 699
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM25
timestamp 1699295625
transform 1 0 8118 0 1 699
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM26
timestamp 1699295625
transform 1 0 8734 0 1 699
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM27
timestamp 1699295625
transform 1 0 8532 0 1 -1444
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM28
timestamp 1699295625
transform 1 0 7976 0 1 -1444
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM29
timestamp 1699295625
transform 1 0 7420 0 1 -1444
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM30
timestamp 1699295625
transform 1 0 6864 0 1 -1444
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM31
timestamp 1699295625
transform 1 0 10582 0 1 21
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM32
timestamp 1699295625
transform 1 0 10200 0 1 -844
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM33
timestamp 1699295625
transform 1 0 5752 0 1 -846
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM34
timestamp 1699295625
transform 1 0 6886 0 1 21
box -308 -339 308 339
use sky130_fd_pr__nfet_01v8_L7BSKG  XM35
timestamp 1699295625
transform 1 0 14755 0 1 439
box -211 -221 211 221
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM36
timestamp 1699295625
transform 1 0 6864 0 1 -844
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM37
timestamp 1699295625
transform 1 0 11198 0 1 21
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM38
timestamp 1699295625
transform 1 0 10756 0 1 -844
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM39
timestamp 1699295625
transform 1 0 10582 0 1 699
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM40
timestamp 1699295625
transform 1 0 11198 0 1 699
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM41
timestamp 1699295625
transform 1 0 10756 0 1 -1444
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM42
timestamp 1699295625
transform 1 0 10200 0 1 -1444
box -278 -300 278 300
<< labels >>
flabel metal2 4388 2027 4588 4021 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal2 4388 -4606 4588 -2612 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 16430 -2040 16630 -1283 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
flabel metal2 16430 -888 16630 -688 0 FreeSans 256 0 0 0 ena
port 4 nsew
flabel metal1 16430 690 16630 1447 0 FreeSans 256 0 0 0 dvss
port 2 nsew
flabel metal2 16430 -44 16630 156 0 FreeSans 256 0 0 0 dout
port 5 nsew
<< end >>
