magic
tech sky130A
magscale 1 2
timestamp 1699112996
<< error_p >>
rect -29 -57 29 -51
rect -29 -91 -17 -57
rect -29 -97 29 -91
<< pwell >>
rect -211 -229 211 229
<< nmos >>
rect -15 -19 15 81
<< ndiff >>
rect -73 69 -15 81
rect -73 -7 -61 69
rect -27 -7 -15 69
rect -73 -19 -15 -7
rect 15 69 73 81
rect 15 -7 27 69
rect 61 -7 73 69
rect 15 -19 73 -7
<< ndiffc >>
rect -61 -7 -27 69
rect 27 -7 61 69
<< psubdiff >>
rect -175 159 -79 193
rect 79 159 175 193
rect -175 97 -141 159
rect 141 97 175 159
rect -175 -159 -141 -97
rect 141 -159 175 -97
rect -175 -193 -79 -159
rect 79 -193 175 -159
<< psubdiffcont >>
rect -79 159 79 193
rect -175 -97 -141 97
rect 141 -97 175 97
rect -79 -193 79 -159
<< poly >>
rect -15 81 15 107
rect -15 -41 15 -19
rect -33 -57 33 -41
rect -33 -91 -17 -57
rect 17 -91 33 -57
rect -33 -107 33 -91
<< polycont >>
rect -17 -91 17 -57
<< locali >>
rect -175 159 -79 193
rect 79 159 175 193
rect -175 97 -141 159
rect 141 97 175 159
rect -61 69 -27 85
rect -61 -23 -27 -7
rect 27 69 61 85
rect 27 -23 61 -7
rect -33 -91 -17 -57
rect 17 -91 33 -57
rect -175 -159 -141 -97
rect 141 -159 175 -97
rect -175 -193 -79 -159
rect 79 -193 175 -159
<< viali >>
rect -61 -7 -27 69
rect 27 -7 61 69
rect -17 -91 17 -57
<< metal1 >>
rect -67 69 -21 81
rect -67 -7 -61 69
rect -27 -7 -21 69
rect -67 -19 -21 -7
rect 21 69 67 81
rect 21 -7 27 69
rect 61 -7 67 69
rect 21 -19 67 -7
rect -29 -57 29 -51
rect -29 -91 -17 -57
rect 17 -91 29 -57
rect -29 -97 29 -91
<< properties >>
string FIXED_BBOX -158 -176 158 176
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
